PK
     ���Zf��g  �g     cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_0":["pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_20"],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_0":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_1":["pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_17"],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_1":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_2":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_2":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_3":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_3":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_4":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_4":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_5":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_5":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_6":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_6":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_7":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_7":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_8":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_8":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_9":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_9":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_10":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_10":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_11":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_11":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_12":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_12":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_13":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_13":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_14":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_14":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_15":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_15":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_16":[],"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_16":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_0":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_1":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_2":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_3":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_4":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_5":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_6":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_7":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_8":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_9":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_10":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_11":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_12":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_13":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_14":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_15":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_16":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_17":["pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_1"],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_18":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_19":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_20":["pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_0"],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_21":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_22":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_23":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_24":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_25":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_26":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_27":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_28":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_29":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_30":[],"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_31":[],"pin-type-component_902067f8-c651-4216-8af9-ec7a733dc9d6_0":[],"pin-type-component_902067f8-c651-4216-8af9-ec7a733dc9d6_1":[]},"pin_to_color":{"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_0":"#FFE502","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_0":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_1":"#0E4CA1","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_1":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_2":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_2":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_3":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_3":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_4":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_4":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_5":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_5":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_6":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_6":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_7":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_7":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_8":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_8":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_9":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_9":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_10":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_10":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_11":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_11":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_12":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_12":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_13":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_13":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_14":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_14":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_15":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_15":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_16":"#000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_16":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_0":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_1":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_2":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_3":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_4":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_5":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_6":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_7":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_8":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_9":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_10":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_11":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_12":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_13":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_14":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_15":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_16":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_17":"#0E4CA1","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_18":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_19":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_20":"#FFE502","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_21":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_22":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_23":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_24":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_25":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_26":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_27":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_28":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_29":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_30":"#000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_31":"#000000","pin-type-component_902067f8-c651-4216-8af9-ec7a733dc9d6_0":"#000000","pin-type-component_902067f8-c651-4216-8af9-ec7a733dc9d6_1":"#000000"},"pin_to_state":{"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_0":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_0":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_1":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_1":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_2":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_2":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_3":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_3":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_4":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_4":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_5":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_5":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_6":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_6":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_7":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_7":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_8":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_8":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_9":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_9":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_10":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_10":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_11":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_11":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_12":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_12":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_13":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_13":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_14":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_14":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_15":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_15":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_16":"neutral","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_16":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_0":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_1":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_2":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_3":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_4":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_5":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_6":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_7":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_8":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_9":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_10":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_11":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_12":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_13":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_14":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_15":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_16":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_17":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_18":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_19":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_20":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_21":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_22":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_23":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_24":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_25":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_26":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_27":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_28":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_29":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_30":"neutral","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_31":"neutral","pin-type-component_902067f8-c651-4216-8af9-ec7a733dc9d6_0":"neutral","pin-type-component_902067f8-c651-4216-8af9-ec7a733dc9d6_1":"neutral"},"next_color_idx":4,"wires_placed_in_order":[["pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_0","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_17"],["pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_3","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_20"],["pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_1","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_17"],["pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_0","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_20"]],"wires_removed_and_placed_in_order":[[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_0","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_17"]]],[[],[["pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_3","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_20"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[["pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_0","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_17"]],[]],[[],[["pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_1","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_17"]]],[[["pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_3","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_20"]],[]],[[],[["pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_0","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_20"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_0":"0000000000000001","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_0":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_1":"0000000000000000","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_1":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_2":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_2":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_3":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_3":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_4":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_4":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_5":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_5":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_6":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_6":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_7":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_7":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_8":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_8":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_9":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_9":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_10":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_10":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_11":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_11":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_12":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_12":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_13":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_13":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_14":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_14":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_15":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_15":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_16":"_","pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_1_16":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_0":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_1":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_2":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_3":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_4":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_5":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_6":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_7":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_8":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_9":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_10":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_11":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_12":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_13":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_14":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_15":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_16":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_17":"0000000000000000","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_18":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_19":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_20":"0000000000000001","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_21":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_22":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_23":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_24":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_25":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_26":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_27":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_28":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_29":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_30":"_","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_31":"_","pin-type-component_902067f8-c651-4216-8af9-ec7a733dc9d6_0":"_","pin-type-component_902067f8-c651-4216-8af9-ec7a733dc9d6_1":"_"},"component_id_to_pins":{"2baf8853-ec01-4f6d-81e3-1b674647738d":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30","31"],"902067f8-c651-4216-8af9-ec7a733dc9d6":["0","1"]},"uid_to_net":{"_":[],"0000000000000000":["pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_1","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_17"],"0000000000000001":["pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_0","pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_20"]},"uid_to_text_label":{"0000000000000000":"Net 0","0000000000000001":"Net 1"},"all_breadboard_info_list":["a4108921-5475-4559-99bb-2167379b2515_17_2_False_670_144.99999999999997_up"],"breadboard_info_list":["a4108921-5475-4559-99bb-2167379b2515_17_2_False_670_144.99999999999997_up"],"componentsData":[{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"A000066","displayFormat":"input","showOnComp":false,"isVisibleToUser":false},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"Arduino","displayFormat":"input","showOnComp":false,"isVisibleToUser":false}},"position":[1086.25,237.5],"typeId":"23db5403-7550-740c-a02b-8b3755757442","componentVersion":1,"instanceId":"2baf8853-ec01-4f6d-81e3-1b674647738d","orientation":"up","circleData":[[1067.5,380],[1082.5,380],[1097.5,380],[1112.5,380],[1127.5,380],[1142.5,380],[1157.5,380],[1172.5,380],[1202.5,380],[1217.5,380],[1232.5,380],[1247.5,380],[1262.5,380],[1277.5,380],[1013.5,95],[1028.5,95],[1043.5,95],[1058.5,95],[1073.5,95],[1088.5,95],[1103.5,95],[1118.5,95],[1133.5,95],[1148.5,95],[1172.5,95],[1187.5,95],[1202.5,95],[1217.5,95],[1232.5,95],[1247.5,95],[1262.5,95],[1277.5,95]],"code":"511,folder,{\"name\":\"sketch\",\"id\":\"e14b3f02-82fe-4fd4-a29d-28c8fc417fef\",\"explorerHtmlId\":\"a8d4f925-7fe4-4c0f-907b-db4a529ea5f3\",\"nameHtmlId\":\"7a49556c-c115-49a1-9206-1a0d4bb8661e\",\"nameInputHtmlId\":\"964988ae-3bae-4cfc-82f2-b6a56b1c9b44\",\"explorerChildHtmlId\":\"91017a22-582e-441e-9168-e0a4f4ec0713\",\"explorerCarrotOpenHtmlId\":\"a8d32b82-4dd1-451c-b8f6-6642612de027\",\"explorerCarrotClosedHtmlId\":\"b1eaeb58-ba64-4031-8ac0-9de41b2d23bc\",\"arduinoBoardFqbn\":\"arduino:avr:uno\",\"arduinoBoardName\":\"\",\"arduinoPortAddress\":\"\"},2,428,file,{\"name\":\"sketch.ino\",\"id\":\"6d553db8-0c4f-49d6-ab17-1d572b0b3bf0\",\"explorerHtmlId\":\"1a291a64-8b39-4a3c-8044-baab2a889f95\",\"nameHtmlId\":\"972543ca-ef34-4c11-b20d-33f6a2fdf7e4\",\"nameInputHtmlId\":\"c230cb82-9ba5-469a-b9ce-29948beaba9d\",\"code\":\"int sound_pin = 11;\\n\\nvoid setup() {\\n    pinMode(sound_pin, OUTPUT);\\n}\\n\\nvoid loop() {\\n    tone(sound_pin, 600, 500);\\n    delay(500);\\n    noTone(sound_pin);\\n    delay(500);\\n}\"},0,252,file,{\"name\":\"documentation.txt\",\"id\":\"8ea0f580-14c2-4799-a918-783e64f4a4c5\",\"explorerHtmlId\":\"c6659e69-dc69-4265-803e-0f78f0733544\",\"nameHtmlId\":\"b03121d6-4728-45b8-bbd3-69bf341d0e76\",\"nameInputHtmlId\":\"42a3ee1c-c5b2-4447-a10c-0f5f644bc2cf\",\"code\":\"\"},0,","codeLabelPosition":[1086.25,80],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mode":{"version":2,"id":"mode","label":"Mode","description":"Buzzer operation mode: \"smooth\" or \"accurate\". Smooth sounds better and is good for simple, single-frequency tones. Accurate mode is better for complex sounds and will accurately play the sound you feed it, but it may add audible click noises.","units":"","type":"string","value":"smooth","displayFormat":"dropdown","options":[{"label":"Smooth","value":"smooth"},{"label":"Accurate","value":"accurate"}],"showOnComp":false,"isVisibleToUser":true},"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"1739","displayFormat":"input","showOnComp":false,"isVisibleToUser":false},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"Adafruit Industries","displayFormat":"input","showOnComp":false,"isVisibleToUser":false}},"position":[574.8475825,162.4985779999999],"typeId":"d4d25393-b9c5-8b08-c34b-13713d35a739","componentVersion":4,"instanceId":"902067f8-c651-4216-8af9-ec7a733dc9d6","orientation":"left","circleData":[[662.5,169.99999999999994],[662.5,154.93473949999992]],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"70.00000","left":"504.37008","width":"813.12992","height":"335.00000","x":"504.37008","y":"70.00000"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#0E4CA1\",\"startPinId\":\"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_1\",\"endPinId\":\"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_17\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_a4108921-5475-4559-99bb-2167379b2515_0_1_4\",\"rawEndPinId\":\"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_17\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"692.5000000000_170.0000000000\\\",\\\"692.5000000000_65.0000000000\\\",\\\"1058.5000000000_65.0000000000\\\",\\\"1058.5000000000_95.0000000000\\\"]}\"}","{\"color\":\"#FFE502\",\"startPinId\":\"pin-type-breadboard_a4108921-5475-4559-99bb-2167379b2515_0_0\",\"endPinId\":\"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_20\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_a4108921-5475-4559-99bb-2167379b2515_0_0_3\",\"rawEndPinId\":\"pin-type-component_2baf8853-ec01-4f6d-81e3-1b674647738d_20\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"677.5000000000_155.0000000000\\\",\\\"677.5000000000_222.5000000000\\\",\\\"1103.5000000000_222.5000000000\\\",\\\"1103.5000000000_95.0000000000\\\"]}\"}"],"projectDescription":""}PK
     ���Z               jsons/PK
     ���Z^8�H  H     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"Arduino UNO","category":["Microcontroller"],"userDefined":false,"id":"23db5403-7550-740c-a02b-8b3755757442","subtypeDescription":"","subtypePic":"0b351edc-7875-4477-b820-546ce15be531.png","fqbn":"arduino:avr:uno","pinInfo":{"numDisplayCols":"29.5","numDisplayRows":"21","pins":[{"uniquePinIdString":"0","positionMil":"1350,100","isAnchorPin":true,"label":"UNUSED"},{"uniquePinIdString":"1","positionMil":"1450,100","isAnchorPin":false,"label":"IOREF"},{"uniquePinIdString":"2","positionMil":"1550,100","isAnchorPin":false,"label":"Reset"},{"uniquePinIdString":"3","positionMil":"1650,100","isAnchorPin":false,"label":"3.3V"},{"uniquePinIdString":"4","positionMil":"1750,100","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"5","positionMil":"1850,100","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"6","positionMil":"1950,100","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"7","positionMil":"2050,100","isAnchorPin":false,"label":"Vin"},{"uniquePinIdString":"8","positionMil":"2250,100","isAnchorPin":false,"label":"A0"},{"uniquePinIdString":"9","positionMil":"2350,100","isAnchorPin":false,"label":"A1"},{"uniquePinIdString":"10","positionMil":"2450,100","isAnchorPin":false,"label":"A2"},{"uniquePinIdString":"11","positionMil":"2550,100","isAnchorPin":false,"label":"A3"},{"uniquePinIdString":"12","positionMil":"2650,100","isAnchorPin":false,"label":"A4"},{"uniquePinIdString":"13","positionMil":"2750,100","isAnchorPin":false,"label":"A5"},{"uniquePinIdString":"14","positionMil":"990,2000","isAnchorPin":false,"label":"SCL"},{"uniquePinIdString":"15","positionMil":"1090,2000","isAnchorPin":false,"label":"SDA"},{"uniquePinIdString":"16","positionMil":"1190,2000","isAnchorPin":false,"label":"AREF"},{"uniquePinIdString":"17","positionMil":"1290,2000","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"18","positionMil":"1390,2000","isAnchorPin":false,"label":"D13"},{"uniquePinIdString":"19","positionMil":"1490,2000","isAnchorPin":false,"label":"D12"},{"uniquePinIdString":"20","positionMil":"1590,2000","isAnchorPin":false,"label":"D11"},{"uniquePinIdString":"21","positionMil":"1690,2000","isAnchorPin":false,"label":"D10"},{"uniquePinIdString":"22","positionMil":"1790,2000","isAnchorPin":false,"label":"D9"},{"uniquePinIdString":"23","positionMil":"1890,2000","isAnchorPin":false,"label":"D8"},{"uniquePinIdString":"24","positionMil":"2050,2000","isAnchorPin":false,"label":"D7"},{"uniquePinIdString":"25","positionMil":"2150,2000","isAnchorPin":false,"label":"D6"},{"uniquePinIdString":"26","positionMil":"2250,2000","isAnchorPin":false,"label":"D5"},{"uniquePinIdString":"27","positionMil":"2350,2000","isAnchorPin":false,"label":"D4"},{"uniquePinIdString":"28","positionMil":"2450,2000","isAnchorPin":false,"label":"D3"},{"uniquePinIdString":"29","positionMil":"2550,2000","isAnchorPin":false,"label":"D2"},{"uniquePinIdString":"30","positionMil":"2650,2000","isAnchorPin":false,"label":"D1"},{"uniquePinIdString":"31","positionMil":"2750,2000","isAnchorPin":false,"label":"D0"}],"pinType":"wired"},"iconPic":"e0155ecf-753f-4e63-a512-9d8bb2c3e0aa.png","properties":[{"type":"string","name":"mpn","value":"A000066","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Arduino","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Piezo Speaker","subtypeDescription":"","id":"d4d25393-b9c5-8b08-c34b-13713d35a739","subtypePic":"b909fea3-6005-4c04-81af-b407c7630414.png","category":["Output"],"userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"494.99052,0.00000","endPositionMil":"494.99052,-114.49945","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"595.42559,0.00000","endPositionMil":"595.42559,-114.49945","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"10.90000","numDisplayRows":"9.39700","pinType":"movable"},"iconPic":"ead4476f-8cca-47ed-b51a-2c979a8b5414.png","properties":[{"type":"string","name":"mpn","value":"1739","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Adafruit Industries","unit":"","showOnComp":false,"userVisible":false,"required":true}],"propertiesV2":[{"version":2,"id":"mode","label":"Mode","description":"Buzzer operation mode: \"smooth\" or \"accurate\". Smooth sounds better and is good for simple, single-frequency tones. Accurate mode is better for complex sounds and will accurately play the sound you feed it, but it may add audible click noises.","units":"","type":"string","value":"smooth","displayFormat":"dropdown","options":[{"label":"Smooth","value":"smooth"},{"label":"Accurate","value":"accurate"}],"showOnComp":false,"isVisibleToUser":true}],"componentVersion":4,"imageLocation":"local_cache"}]}PK
     ���Z               images/PK
     ���ZP��/ǽ  ǽ  /   images/0b351edc-7875-4477-b820-546ce15be531.png�PNG

   IHDR  u  v   ��:   sBIT|d�    IDATx���}tSwz/��$۲0���Mblc0fB��3���@��0�b�!d�qN�bν'�tAgڣ�rf��i��Ճ���M�8�Ms�z��� N�`L�~��-�/��ClE�e[/{k���Y+kY��O��g?���S��ҡ�D�P�C���{HDDDDD�;����_��{�R�=�p����V)v9""""��Ή�:�t(I�R�)xZ�Q��5�cR�GBנP�@��x�1�cR��+o6I���t�|�&�I ����W��ǙM~��<>/(�^h�J""""
O����=�p���`T��F��:ix./M�8�IV�0<<,�0������ ~�}�M�Kb�J�/^:���Q��)��ӣ ]��+���!�L-[�,(q��~cP�Qx��+u>HT�*�GT�K�N�F#�0�����BN�T���@{��c�NQ9*���!�S�=�p�n�DDDDD��abg�{�aR祄W��="""""�G('v�~I�v|b��
[�M�6ן)�B�;JX�&"""�^�N�dRDO�f੅�`�b���y��A�����DF=T*~��"�bb�������_��g}� �L|v;>��f�@�|y`��6��~�PN�JU�Pث�B�GIDDD^B1��^Jx�PI�g9������~�1��y��\oo/���@�Z����80w��Y���G'Q�f
���c��	��0����'�C
���䎈��h�P�:�aLv��0�Ə��8��/�ҡ:m�Ҡ ^��٨���w��cqyX˸�˸�Ըb����q7��
B�b�J��X���Z���qu\e����MRʕP��{`<�}���R�a��A�<�,]�q��G��s"�������m>=?*v�~I��v\���H�����_�W�J�@�g�DDDDA
]1���1!����(F~�r;"""���N���);`W�*���	F~�r���`�#"""

�r�f��0e�tk�f����봯��f �S&&�ݮC�RA�R1.�2.�W,6����O�P ֋�y�q7��I��f��b�`xx `�Za��  � ��������"��<x��:�����e�?�S `||f�FGGKllRSS��!�2.�2��q�b��1:j���H��R*��?���\�e\�<n8`RG����`�Zq���ޅ��?�6�������9Z-���/��#�uB�)�o�<`�P�B�|ǟ_W*�P��D h��q�?>�v�Wg�˸�˸���B��J�9s�tA*\����xu1ʸ�˸��L���������z��c;Vcn������ݻ���|���>�����ݻHNLD�R	����	L���X`������͎/&&�y��]�����BZf&������(�k�Z���?}(��"<����8f}��6��1���F�oV�[���pa�P(`���q�q%�+�@.H]/D�q7�qCYd���fý{���ڊ�`�Ղ�y�H���%&c�}p���� ��#QJE,���0������F���`Q����b����ܩ����)lF��� 7&����q�q7Xq������˸��	���&A[k+�:��א9/��x���`��8J qJ%�J$ƨ`�����������'�=�RRR�z���.�Z��ƕ6c�MPR8.�ZZZ�~�ʕ�D�0c\�e\ƕ�J����;ר�fɒ<Q.D�q72ӟ�|U��Ʉ/._��cu��j��Q����qc
̍�A�J��]��f5z�菡/-EFF�#�"v4�=W#�x�I�ꛦ@�`
�����&�)�e\�e\�X,V�_���~�q7��"��d��_��G���I0wv`��W�1
t11xT���}�O���B{{��1"�ݎ�oa0�K4������:��d�o��a�ڄ�9��&��$�� �T���x�_���＃��nIbE"��� �&�D����(�0��r###�M}=p���`W�A(M�*H���D�u4��?��ݻ��$""""�DLꢘ�f���1|�7��SWWP�����k���gQ6��t��W��!Q4aR��Z[��#;I�� 't�X�ɱ1�{���ٳA������(0��R###�ZW�m"�;�2�r:j��qq���Z���m� !�r�a2�MY"��������(����B�sc����e��F��vxW~�kV눈���|��.
Y,�7��|�C==r�c�����~�vÜV(V��ЫE&uQ���Z�#���N��,N�D�݆�S��J�
�J���@DDD�b�@4��ݥؖ�,�Y��5O�C��`���54`�ܹ�Z���
�����s����{H�'��9?>T��A'Ʊ��ӽ~nll�!�q�qe������u			�˸�BqC�� �L����z����_H�X,�tu ���m0�X��!t~�%��^QJn
@7��C�^�N� @�MY!�q��Ұx�b�~gxxV��7H�q�qŌ+�����;V���Ì˸�+s�P��Q���/��T���/�P<�Q*�Q����,�PB��.N"%��@������D�/!!j��q�q7hqŒ��������{j�:�J�2.�7T1��2��혫���phn���cm]��~'�PB�B�����=��WU(��K/��^�1.�2.����Q����˸�x�P��Qftp�PȾ��LT
��^ht�Uj��h����^:��P(���u�J����.�			���^Mkf\�e\��5�X
E��!)�f*)�2.�70��2C�3�'�J���.���(xZεu��!�*]LLFGG���+�x�v;�2.�2�$qŢT*#���q�\1��211*����ƬT
�G��P���P��/^n
fܹ�*W /r�͆��Q��ĸ�˸���v�,�g\�e���5uDaJ�b&�F�t()X1���P�Jc�����E�ؘ�(�*Y��B��J���nΏ�ؔ�6G!""""q1�#
sBb7�Ǉ$��oʙ����(ېh��j4rcF���,��B�@A�Mِ��������])�x�P�æ(~�����w2�����:�<�������a1.�2.�J�A�<|�rیω���q7��"^9{)��C%1P�	��K��?��Ǽn����+z�իG��~��|y��	Q�-���	Ld/Ď��I����%9n����Ʉ�f~��@���ʡ
�BiP EQD3���,�+uQF����/>Gl|<F����G�v;�͐{aK���1P�Ѿ��'v،C�Û/x���ĩT�
����Qx`Re2�z|u�#h�ڐL���vL���Z�B=�O+�|Z�w쯼��ݎ(lm6�\����

{�(Q(P L�%"""����.�:�ڝ^<��>�R?O��&��		S�#Y����;�?P�v;,6;�=���P�i�Oʩݑ�8N��Z�>��  �ͷq����#"""�hƤ.����M��ۛ^=�؎՘+�ǳ`u�?�-�B�Z7f�#5�		r�h���4��� �Ä �m\���.�2��,��`�Z�����Iu46m�5�������CDD���A�{�i�3����*�P܌���۠��?�{(DS�4jԾ��-��.@��2��I5�v�PV���t�ㅙ�0���/+�'""���J]R'$ ��߃��fHU�6�s�h�j��B4E�~1����� ��q ���#;E���AY�竺=ې�Q��ݏQw���gBbW�gJ�����$�()�%i�����ꛤQ���#�����U4��`	�����I]�Z�y3>�������H�6F�6<U�W�y����6��Q�� P�w�3�[�� �a�ԕ�03�oECKǔ�7u����h����X��3Wd%��$�U��P���V�0[��kB��IΧ$�Ez$͉��B3�zM0�;Ө��ك�O���G�؁�Y}�rпk9�:6?�f4�t�� �9% Z:`�o�}��1���P����(�#'U��7�a8�i�n(5T� �T������R�π�]����Iա��է/OIn�vJ���Caf:*��(�L��A��I]�R'$������e$��b�����2a��j�!q�rV�$�؍ӈ��t�Q�|��4�q��}�^??ntK��J[`�1��[U;a�o��TI�03M�=��.�"�@W�F� �]��8V,q\��t�$/��b�����9�Iա�j�󮼐 U�_���-h�Daf:��lsܬ��.I�FyAJ�fKrq�� ��B3J�`ܽ	m�&�w�|��+�B�!$��bT�_����]��$�%yYh�ډE;O�d���1�p�ؚ<��_��B�]Q���B���)�����s~�m�&g���HҨQ��.˿CR�(ңzG)�zMh���o���AR%�rbR����p��e��Q��`�b�� ,6�J��/�"�����'��^�Ռ��x�I|��Ը��� ��+nt�>���:���˜�i��P�w����[��:��iҜx���L�<�ԫ��:	��s�*]����b�P߈���h�쁡����0�����fA����8Ū�+U�IS���ls\ؾ��(q�V���0l~ʭr"er'�o%�G0`�¸{�:{�>��ӗ/m~J��M8\+w�k~�><-J�$�U�W�����g����U��r$�6!�5�7:���F��)��5l~����`��*�^�S��*�����2�Z���|�#�%��(�����?�	]����ڂ�ؙ'&`��P��͎�+����^%vb��&�3�s����Gб�ȹ��5����h=�t�^��4���gO�	�J��=DI^�ǋ�����VSg���\����k�����f���:{P��%JL)�XP��Ǩh�pT�&�-h��ASg���sRu��v�y��1����vK��-I�vN��:��B3�o�qU�v�#BE�����b)��r;?��\q|��r{�����Ϸ���oEݞm0��$i����9��k
ڍ:�����^�O��o-��(�NH��?z	��7�@F��:����Yl6Xl6<��z}PbF#�+�l��TqgJ�H��wocw�_���6�fck*��=f��4���#p�J'֜T�E}��V���rR�n���z��
����sKĎ+�f/4;�r����V �zMn�[CKrR�S�����dm[E��9�q��b^��A��M0���V-��b��n������3��{1�}0[Q��ǎX{�IV}5�7b`Ă��U(������0[��TeMҨk7E�Ć&u�y�����������I_��yX���{�R��g���J��%vR����I��	�_b�K?F~َ��|���:bO���iHr�<����6���]mA��RwoBCK�V��X��<����C��R��e�����ݛд�nu�;J��ԕ�WjBr��Q�di�#����B3��ls�w���>V�_�;'ޙX�y�?0b�m�p�w0[a�Ќ�T�֯���j�5���0��PV�ܣS*7�a(+F�ي�3W��h)/�s~O�|�B\C� n�;oX	�_��I����Q	��N&�$�I�:*ۓ�/���(_����Hä� 8���j���~�0��+I�q��	&�
<��V�$$ub%���+�kb���5���Q/A�`�xu�t�l5ቶiH�;J���O�i��tęr���	�/��W����3WP^���-�><-�U��T �)�U�v$)��-q0�7��܀�*��.W-�u|�;���*li"�6�7����/4;�f��%VBYx��VT}x�ys	�d7w��\AҜx�t�����K�r�|��g�8���,�ñ�I���ZQ��<�B(܌��j'>����r \$�z�$�3��wl�j̍~�mƥ�%l-7��h���=Q�����0n�#&�Q���	�����{�3u%�=v�44#��[̔�(�FG���#K��ێ�1K��v/X���&i�h{mϔ��+�d��<%u{�9�	�֯Dݵ[nI�q�&$͉w�o�".�m���ׄ�w?F���:���H�`�-�3���>(���C��{��J�4'^�q�$'U7�1�	[P��3j��A����_�
	^�>/�r/l{!��TF,S���3.0��Y�~%��e=�� |�#4u��|6���,�+u�F���5�{��܌k�|Z�s���N�d�f�æV���ǲ?�C�Nn�>���1Y�&<�J��S\MW�4�����d`�"ZBmӐ�F0u{�9���0��n�6g�W9)Z�,�FI^�dӢB�1n����dO8Z:B�
�{������ӽ.�_�lǏ��P����*ؘԑGz=2~�:���q���	�qq�%%�n�atx��a�'<_H��혰�a�c:[|<����d�ȅ�{�T�gm�-���<�8����g�8�)��t��>ga�]�$_DDN����/����S��e�����`�b��4�S������9|s�"�{�C��F������v�Y,Ǹ��ݎ���1O��%6bޢEr�I�R����bb�������_��g}�߿/P+��C51Ԙ�΃�l���-�Y���ʊ�����$R�]7[�Nh�`Jw8��G�4$O�w0M6\�1���(Zp�exj�#���{cc�]|����LR������ہ�۝�u7O�뜺hQH�7�]˳�����s������ΰL�����q�g��{}&��[�M�x	ӳ�O��ݙ�����~��;�q=6�u]�S^���M������R�]7ݴ�$�ڹg��Y�S��q�X��|%U����g��d��w#�N�F~Fηv-f��'��z)��ԑ�ع2��$�Ŝ9j|��9ѹ�g��3l6qo8���0G��Wmw<�������fO��!n�(/ȃa�S���"6��tp�:�.@s�}��|+�!/?#�+� ���j/ݐ<f��'��z)���E����P�Th���x��=��B9?]U����F��U��u�~q��2�&���q��Ձ��w]!6/_��Wc߱��� q]ﾇ���b�'p���o�-y�q��E<��2<�jYT�'�ߋ�[ס��)��kr3 &�U�}]�3�P�w;��q3>��ɋ8x�d㐋R����j��s�O����R�".���_$�E%yYh���l�!eB8����$��q���|k'v�s��B�B��lE͹&�w� ���ηv:�h8O\���Z�G�6����gp���{�9g�'o:aL���:"�($T�=ڂ��J���|�ś�w�I|k���E�yM�7?#mJU�sּQ+I���ϭZ6��-���Lꈈ�����FU�WN��^�y�h�ϸ�$u{� ���,Gv�Źp�s�^
��q-�I4}/jvn��XVr�dSm���2}�պH��ʤ��H&����=�$�;0b	�F�MXrRuAm�ϸ���������}?**�b�êJ���-�[�,jΓh�^�۸��y���Bo�-z����A��8�uݴ�9��m�7��7T0�#�r�� !�}Ͼ�ix0<����q A��i2{�Ed\Wf�Ǥj��DW��+�����\�578��uT#��L���;�F��V-CG�P�.z��<����i��dRMì9ׄ-�\�.��A�h�V� &uDQ����T*��
T*�����װXş��so��I��TJ�`�"\��+H1�]����T	N �����T�����ͷe	y���,xU�h;O���z�v9���0+?8���2��ȩ��F�I]��Y>���Gg��y�wa�\uF]������סP��P�����4�Q��~�l�	���i��$g>z�� ��>���mbv�j�������Nː+n�JҨQ��9�:�TA�F��Mn�ih�@��Ge!�3��q��ͬ���nv�:�:(��z�D��n��d��|\����4�H�v)`RDm�Ch���;��G֜�ٟH>��l�|g@�a����<����<���;���6H Q    IDAT,$͉��}2I����-�v�LҨQ�g�c��ӗ�~f�oD[� rR�Ά*rOդ�s�l6/_��Ϡ��e5�=$����{hl������k{���W�'�v�8y���?�_ock��鏮-��w���Ps�	�cZ��#�:""��`ܽɹI���R��}Թ��� ��O!'U'�vEz����	����J�f�di6�:����N���e�;�1��j>B�>����?(y�h;O�����|4�~t���h����D��:""S��0[QQ�w$y~����(ң��G��K�f��f��0n���t���)z��F�EU$�on�4�h;O���F���PŤ��H���>}�Y6��۳%yY�>sE�΅I���n�lE��+n���"I�F�F͆)�N�bתe0����|#���������o��cDD<L�\\\�^4	�%8���&$Jm.SO�d�03]�ꜧ1L69��9&t��N�:[|?���X�F�,����jl""
&u!*F��J5}�>�(�ʐH�
EP^/Q��>}Y��j*���>�$/K�M�#���N$��ߢ��-ؼ|1��fmz����i��1Q�aR���P��������oJg6��9o|�	��A$�6��@ݵ[�*]��������T�_��<T�����&׺�a��ŲĖ�)ɇI]����\�+}��K]}���F��0�o�Z�aE��^�O_���%yY0^hv&�9)ZG�ˇ���y3�=���  K��L��A�(�tDD�I]���i�_���AsHT���j�JT�_9�c��FѧdV�����AT�a(+v�Y[�	��Fne �5���JN��An� ��\���D�]�����:"� 0[=�U�����-��ڂ�T�s���^��Id��f%��?�ڿ���IQDbRGD$���#^=/'U��i;ö����k�4F��i�(�]�����O��HCVr"���s]E�.���řIQ*/�C��%�f%\���3�  �]�"�u/l�MD��03Ezf�;g�q�zM����K��E��<wo���-0�7�M�2�ބ��[R}��w�֯DE�9��o�s�ٱF��n���S��L&��i{m��}�\5u�x]� 
G����d.'U��^���p�]�Q��w�àe{�9���^���Y{�#��uO@�Q56E'9���"=�w�:f��N9~I^e�(/ȋ��I&u��̕)�f�ø{��lC�ύS�����^�=�۳9)ZN|���P��U;QR}d�4.o�9��۟�^ۃ�^SD~�&�Z���qpL�du.���V�;�	n}�6���֮�%u}����)YbQ��+��(�;�a�a+���,��ن��+#�bǤ.J4u����T�(u|��8�K�P����O�]l
���v::�M��}�$/�Q�+�C�F�'͉w��Ä.��^���K7�.6E9��$�������M�=H�p�Pä.��8Od��<M�l��Aҟ����#�"I5��ls�l9}u�n9+ܳMY&""
Ur%Wf+�Vf��xS4I�v4 ���L�HN� ���p��Q�++FN�M�=0^hs�DQ������>IDDaN���x�U�W"'E����M�f^����K�ύ4L�DyA*����������﹖��VT��1eŨ(� �w����-�>}��<��M��.f딵tD�"��FE��y��Q
CY1�Qؓ+�2�7b`����Փ��-0��4"�8`R��֯D���S��D��QJSg��>�$�U����Q;�U�Q���)���g��0^hFaf:J�]e�VʊQw���QX�3��>s�g� 'U��usĂ�Ξo�"i���1��@��/sRu0�ބ$�zʖ�0[�1�><�ܾ�zG);V�������H�Ҡ�H���+��ك�w?���DD6�M����t�������$��?���+80��p���?,Gݞm+iު۳����LV���l��w?"ѳ�O��ݙυ{��ۯ�7w7Hꮶ��j��
^^����t&uDDv�K�b]3&i�0��03U��x̊"��Y$΂aR烵smXk��ܤ���VǨ#�N[�ɱ��mU�n�;۰{��!̝fBRRt��Q᫶;~�����f�˸20[�w:���7��]1f�U��B�_V�m�%$|Ez4�t����y��I��~�j��Z�q�Q�R���������!��KN��U�(EN����MҨ���P��Q��N����*F���>���	���䬘U���hܷ��ݛ`��r$q�W:�Y�E"&u^���~�slԺD�q����Ά&��#���%�F���Z���	8���T��圮�%��2s�����7w{�S(����|#w�L��4�;�W�zM(�(Z:D�j��yA�T�(��Qw�I���''P�~<ܲ�[�N	d��: """
?rW�\��������C��l&uDDDDDDޒ�b�:�L�V�(u&���� �oq���*fR��Q���h��A�ύ0^hƀي�w?v.Aj�ډ�"�dc�+uDQ���Hиw|�^���C�0.�$�3a C}�ǥ?���)��;J1`�F�>u��E��{C�J9���:(X�	s������&G�l�lE��Gg�� L��ԭ�X�#�R�{�`��ݮ��9K-D�o;��H���df+�O_�r�iܽ	%K��4+/�CE�%yY��ꮶ����.Ԯ�_�~�[�jO\�XW�(����(�c��U;a�oDCK�v:��=����F4u��j�JT���������nݼ���
�I����ԡ;'U���?���᪢H��<Y����b&��+��BҜx��MҨ��Q�/�0�#�R�rL�;U���h���PyA��BN�n�}d�d�P��h��m��9m#����^���i��䡩�Ǒ$�T�0�����6>O���7��{
�M�=HҨQ򰃢�di6�V��e�%u���h�5����L��MN��W,���q�¾�Ez��&��\���i�#T�f��૜T��>��(���sw��E��K��/����dUw�����H�r%(�LwV�\-�B���U���0-�P��hn�R��P��&A4��9�:�䡡�f���"�����)�7&'����4կ� o��#�g����-��܎���&7s�sv=��1�����%i��
�l���&W�;J���s��p͞��>���
�4�H�ހ�:""""��]mA�槜2O*��h�왶�2y/Z	chh�pTU&W�Z��2�q�a���,�v&�B�Vw�e��?�ꐓ�CÉOݎ��ҁ�<f�;�ϭ>s�y��wor����Kv��{�C (�<�j[�p�\�[ ϯz��O��b��Z'���t�i�m�&��ن�=�7$�OnL�"Шz4#�݇e"&V���sS��>�jb,�q������3c��$/u�nI:�
&L��vE�Y��Φ�H��؅����4n��U�
3��p��m�eCKJ�]�Uw��m
f��%�W�������2%U�|1��q8x�"���]O.��Gq��.��e�}��g�CG�Z��x>Ea�\[ߠ�1�.�L���+&uD��e�x��$���ĳ�p;� ��w^�,���EX���Ci�j\""�ʹ�+�C�^O����zf�_�ufBu��f;�֯DyA^@S���{la_�~%�֯t{��j�]�Ȧ�geM�
UɆ�gϵ7YCK��rVq��®���Qs�	 P{�j/����L�]W���;�]���'��|�Y�Z�b�W	��B�䛁W���	���(b}���˪N���A��;/��  ���������5.���K|��t�,y��r6Ez���9s�ʖ7rRuHҨ=&��L��Օ�e�-E����}����n��L7ƺ�-0l~
���0[��2��j��
�d�[;q�uj���}'�㍀`��}m��<�s��E2&uDL�krB����`$vL�HJ9)Zgh�!L1�JI^rRu�H�Mi,�4'~��,ꮶ�03I��4N�6�9���칾�%���.���S �����E8���:��ΔXI��1�#")��9�|�0M�x�ٱmA�S!gC[�	�~����f��$5m������kKա���?{��s����j�w�pt��$����*iN���n�ȑ�y����1a��H�����r !!a,!!!V��^zD?2fW���#���?|D�1�;����7��N�fK褊�Mb%EbǄ���TQ�G���0^h������C}#��7�:3�9m1'U��Ι��~_LO׈E��:��K@M;����w���vT��������E�>e�	d���������P(Rl6[�7�x�b���h4���[
 q
;  �_(�a�4h4J ��Ð���x��i�YG:Ψz�\V����N���n闟�������ݛ���g�J��B�W	S��+h�t44��9���2eSs_�����U.��l��p�d��:]zJRZ:`(+�j�_ݵ[���t
3�e�|���G�
�X[z�+�O���6��^�����INN����Wm�
7�Lꈈ�䒤Q��/+P��Ѩ���E��N�JK�3���,��r%"""��!l�0ymI��������������I:Ez��):peE��{
�f&tQ��:"""""�0�JQ��N�";Y+�0�����z�=�"l�s&uDDQ,?#�{�C'�P�������>�j>���.f��#J�|�0Fu:�l�)���f��A�j_������>cn]��#���hX�#�pm��A[�i����T�sASg�c�Ym�+��(/�s�Z����f��n���z0`����e��'i�0��mJ[w��������&��z�8+uDDU���c߱�rCTLꈢ��x5�t���/��S���0��03�~�|�𸡾�ou>nܽ	�ݛP�QO�e�o��
��Iա��� ��=� 8:�5u� 'U��M��a9J��` ��F�������Z��#"���5uD�rRu��Q���� ��\AҜxT�_��k�����U0^h���U��1�2�Q�~�W퓫�\AyA��P��i��03U�FSg ���C}#��l��A��7���A��ADDD~bRGe�֯D�F��ӗ=�|��I5�4j�z^�Zx��>�o�5�03��騻ڂ$����:�4'ާcE#&uDQ�$/f+Z:<�|�l������-(��Bݞmh��P�,'U���Y��03 �������LꈢLҜx�X|���<����F)��b���&)3%h���z�I��xEz������IDDD��Ѭ�VG�w?vLߜ��Y�~�Ǧ(��bʊ����T�3�ބ�Tݔ�~DDDD��:�(30b	h�����Q^��槜�T\;UΖ�yb(+FyA�����?"""�h'߮�D$��k���Q��77YyA�s����+1�7?r�ss;��/4;��4;�qwoB����x�c�}��hfLꈢL���0[QU����'o.4T)/���|��I��v��S�����?@��l�TaBGDDD�#N�$�2f+�><���{�6��SeŨZ�-Ω�M�=�>sŹ����9Ͳj�JT���EN�ι�x��G9咢Nv���Zd�$�m �67�c�\�e2[q��>���k_A�F���4�g̃N����A|��=9��u��:�(Tw�%�&GW���xSg��'��h�5�� m��q>����H��RYQ�G�F�8��8\�Y���~�(�g��L�ks3�� ����_��`ڟ5�v�\k'�o�z�=��*�F�|���f"+9q��)���i�2��8w��[�"�=��������BZF���'��t�,š�Өa��#��_]����4Ծ�Yɉhl�¾cgq��ޔ�w��d�bד˰c������w���[��6>o�k¾cg �6���uO  j/}�|�u���~��'/N;v�F��[��U���?�'/8��؂����®w��z�=d�hQ��)�O�Z�)X��~#b�J��V�|���������O�?��R�@���_��ɏ��DRQ��Ԕ(��3r !!�k�N�P���~�t7�r�(�}�5j�,r{lB��X�bUP)��o�u|jK+���bhb|O[>~���H��u�(��Κ��k�2���V�w�ηvJCj��\�-�\l^�X��w������5Ed�L���[׹%X�V-Á��ܞ����q����P�q�����p�'/�%э�](�����E�s���7p��E\��
�c<y��oLy|�����}�+�q{|��  ��������_!?c�Ǳ��c���n�����7��s��9��"��o���-n�TG���δ�����
���a��_���]n1�q�o~�L<;�����Y�7G��e���/)f��X�#""�'����p{,sI.�sf��x-!6�w����o&�P�%�ZŐ�6>ϭZ6�z�t5*�b�'$KxYɉxqm!^\[����8|x���ӨQ�s��=��������Q:n�L>W�s`Mn��&;y�X�1m�|k��Ǘdz��c ���X� ��؅�ɳ�G�5��Sn���k���@JB<�-��X,w^*�O��ޫ(Ê�#��>&uDD��AF|U� ������^��B��~��I�t��q��8��i���9�$�8f�d�}�<~v�o,
�ؕ0��d�����p������xs딤�d��d�N���*�k�s���8�ډA˨������?5q9���qJ�[���}�㞎8�E��V�c��}oʴda<��p�鷍�]n�����Z&�6�}J��쭎)cl�?�-��)�g'k����޹�N�tR")��lْ�P(*�@\\�)>>>I����}� �-�r�HU�W�_��?�el���}�G�M�&���%A�Pa|�
�Ō����A��>� �`��c�{�F�W���f�~�v<S����Á:F�?xl!��q�����_�!p$��/�������O��{�!��dMn&�� u�
:���B�~��wܞ�x���"I�ƪ��`�2��?:�������7���Y�����͆�w7���|k6<��F���.�?E��.}������څ�N�gh���X�$�[����;�L����:ׄ�'/:�ҝ�:}׻ﻍ���˨�|�ۿ�8�K���;�S����|�|kηv��>��-:�����_��?���������9�������}/t=C#h�@Y�b(
��@�q���.����Y�P(�34�m_�F�5�*�����q��&H)Z���t�����?����#.��Q��:�dU�W�PV��fﮞH�\gw{,1)���n�����I�Z@��a^�b�'L��;_��2�r�G��	SߤZ&���F�S�5w��HC���g̓%�7��%����۸zʚ2!i���63!�6g����MY;(�ף��5uDDRF'�KY�R��Xb����p��-$ν���ˠP�_��K~F��n�m��/6/_��?y�GN����D$�.��Wv��MGX��ӨQ{�\��ų���n��4�pg2[�$k�SovonŮ'���U� ޻�?+7'""�R�e#!1s��	 �զaђ����t\�R1���8�Ņ~b#�]O.ùW���N����{e�ٹa�'� ;E���
��N �G'u^�Cv���݀��Dh�����B���x�e��[皘 ������>���.��5���m�s���L�$
+uDD䗌��ߊo:�����FO����ڧ���V-s�W�dS����n�͋k����uʪ��[��(��ȹ���}�κ}>�nj��]�ۏPhb�����6���`6[1<t�c#r'(�=��3���O^�8],P�k�^EY�&t�����r��v�R��HCv��c2y<D����<u����'��X�#"��d-�.���u�:t����=$�H��]���e�}��kr8��J񼷗?��q�߻e�?�uk��!�{d2[q�ս5���,L�B�-�    IDAT�Q#?c�3�DM���P_�]Ҫ�������{���P޿|��9�2��^���������?CaSw6�!10�#""�`||f`�L`��M����3f(�\[(j�r���o��ý������5��آ_�2�d�J��N�.�׻��K7P����_�b�G��y�ٹ��9�f�k�2�=՞[�Ǜo#��oI��Wy�*�����\���Jvq�ܺ��s"0�#""�%$$  t:Gu�61�ί?C�|xL�l���mA����8 B���A�^���.}�S�⪣�_���/߀6>{�=�]��T�4��iԨ��.�vR�G��|{������qp�:Iײy�0�g��N�$���4����I�F������jo¼�Q�5)��a���m `��)F�)ڀ�E����ɋ�iWb����ɋ8x�"^\[��W�=�0�Į�bK�	����[��ֹ&<�j�o\�wr���B�k�,�:�b���'l*��1k'u�l���}�7<������{���%v\cG�bRGDDS(Uq��O��wU1j<�Y�{�����;�Q١��nj������lE͹&<yQ�QM�hm����k�:�?�]��nS}e2[q��E�6�Ry��c*��uO���B��X��=�6(�i�صj��sq�������w�\��qn]���f߱����t�cp$%�T,'�^{��hS�3�ܶ��vL3Y�����
g�B\�o��A�(j/}���8���#�pp�:d%'���7�wg?þ���{�*|��%""�hS�C��sal\<2�W  ���a}��v&�h�e��B��������~O!�Ǡe������V�<�����6>5;7x�$Ц(�ͭ�<r
��Q���+��y���[|�lj��pp�:���ܺ���.���oL����in窘�b���~}&�^1�x�mQ*�:�:��	�����	{���O^D͹&����7�:߇5��h|e��gϯzܯs���4 "� ��b�͏<�W����q�����ohԌ���qv��C��6%���KG�Qc�������K7������йjl�7j���Ϙ�ڊ-3>'��1B��yc}P:W��]���;~U�6/��)�a$l�1�����E�L*���+�� �۸�����"d�:��zq�I����J��0��Q���z��;��>�l������ߙ�L��G��;�T�o\�״�}��e*�l-��R�+~vv=�{� t��4�mד��n��7�]��hvٚ@.��Q���{}�?�u�(��k��Jr�E��W����bo��Ϙ�׺T]|�$�������3WP}�J���f��ɉ��I]��N��E?֥U9%z��@������ZC�1�c���~��z�=��(�!�;��.���f%'bד�^����'8���?G���x�m�+�bp������o8��:�2;E�5�����=V��Y�z�\�۱�����:""�Iv�q���ҍ�K�B����Pvx׻�!?#�{��U�ńN0h�.�q�Wn�ij���E~'ukr3�������T��P�,����uX�F�,�����޴9��m�;vv�ϡ�o�}�f&kr3Q�s��ݞ�˺T���nKͯ�&wLf+�:�aMnfT�8��#""�d�'|z���N�� �7>x�_	�p�*l�i	����>�إ4+9ѯ�ukr3q���۸�6��?���z�x5Á>c��]Z�Ө�ݢd�����^�[;��Z�S���߇�(�[;q��E�X�����v�|�_�ŵuaH��F9�2�#""r���e>%.Bӏp���S~��g�õ���k/:���[ס�r�����1<����)����^qͤi{��8����f�9���Em[�y�~����_7=Lf+�j>�ؽ����)Z�)���8���[o�|��H�����c���ɋ�u��G�SA[�c2[E�н�p{	O����q:�&蛗/�����]+�pv��gn����I���ǣ�S�����y�K��S�6Q	Or$vLꈈ��i�3n<<Y{�`Ht��Še�GNy����f��e�C>_���?g ��������>�o�t�pt��k��E��!f�)����yڭ'&��c���V-�Zw��ޔ��q:��<���1�#""zhMn�O��bP���%�2���ِض�N^����VwMf+�s��yc=�7�c���'١�Se���uAٻ�S�x������K7<V�}�Z[V��������N�&�n��`&vLꈈ�Z����}�!���'>���)�P�ꍎ�!���r3`ד���k{���#ܺ.��� BE�}����D��)��L�;e-ݠeT�
��)� ����{��&�O^Ĺ[�x~�㨯��J&I#X��:""��|�8��<�����s&�}����{>�/��8���4j�=鲒��F}s+NL�����P�N��n��7��^!��p3#+9ѧ�)e�\غιf�����7�!q#�cRGDD��/�߻�#	�}�>�qJ���n�''>�������OIK�6¨<2�<�n�1x�as\�u�&�����Og����2��Rh�:����DDD�|�=���A�׋��n�&����Lh����۞�^���֮���7�M~F��]=Ϸvz=�-;y�J���Nt��mV}��-"��lŁ��.�/���XG�醍��Wx�xs�xޜO7�K��{��a���*�>6�:"""������rm��E���7����h����ـ*%�u��V��͹W���g����+Q8���uR�671��]���﯆.^�s7��V5皰E��b�*������ۢ�5�tS��H��4��S����8�p��/o�k
�6$$=�;N�$""��)Oӹ�g�N���ߓ�/��r���ـ�]J���{l).�u5�u����Vv6�c��+)�����K٠��/�}+��@V�܈M��)�e(�I1�I|����w���x�N�ӹ����M#�2}.�W>�}W���u�����"B{���je0�����J]�ߚ���sq��]���lG�{Q�&2$�;&uDDD>2Y"sO����~U0"uj�/�G�ur�ٻ������y�X����5�b�]�I��k=}�&o�0��[�9G'i�����:"""r�Te����Q��Gܧac�P6�&�/�y)����1�#"""')׶E�Ó��5�vEl��W׻��I�X{�I�EJ���N�׏"���:"""��s��\�ʛ���ͭX�s#�����BY�GAY�8p�":�ݛ��1��S%y�[����]��8��m4�v���7�T2)���qK"""�g���������� �"l��c�_��&7��/��0�{����u�ZG�д��}o�Y''�J~F��s�Ө�����-&3���<r
�+�q>&��uR���[�0Y��o���F�] �0�#""�o��z��Г��V����Zq��zr�߿_�s���������4j|�ڞ���_�z�����WQ��󾍫a2[�*a����N���66/_�|,н���F�씩7|i��Өq�'/8�4��������E	;N�$""�o�n"m��6>5�6�M�Qc������ƛ�F�^_��y�`&;yj��E����|�V9�vs н��F)v�.X�a��/۠T�-t떩Ϙ�]����B�ǟ��Lꈈ� �6���H�Ey(�ٹA��ʵ�(�db�2��ٟ���^T�<%��C�r+'�ي}�>q{,н�<M���ٻ���;��H���e!"8�Xp�d0�f�T�2"����=A�dfrj5�����`������cMrƐ��(g-r	V0Nl.��E�`ld���ڒ��R_��;�����[?���r�~��<�H����<�'Q�wK�_P!ъ6��  �"�bf�y�g������+�,��mј�#X+y������ӽ:`Ц��X�t��e,�^D���'��x��We4��Eya���F�;9c���P�/��h�� �+����;k�~�"��Ƶz���*��灻�g*<r��:?ҭ	��P�7��;^xY�O�;��������|v��dT��<sf<{�S,����7|�p�$;�����=�Ԗh��Ǵ��c������"v�:  �8�L3O5�)+�k��BvݺV�xP^F�v�yh������*~�a=s�����zC>�Gό*���3򔌑:i*ܼ��3�źw�ۧυ����|5��=q����w�=֕�ЁǶ�ÿo�-�Wh��"
v�:  ����}�����0Wm���Ѝ��<pg�ih�Z��f�7��ĝ_��o�ᕤ'f��3 X�蝹f+/#ݐѺ���z��>l����9k=Z�{ׅWO���
��.p"M}mF3���c�C�?��zC����p�`G� ���'��ւ���I^F�<�=��N��h��%���myံ��i�?[^8`�3�����Ϳ�k̺�x��4'�>�A�g�q�'"�jj��oה��4�y��9}oe͠ue+�Nen�<�(�����k�`G� `�h@�����*��{]o���L�ڞ0&�u:���sa�9=m�C�Dx{�F�9����!��}�v����F�֕��3�6�,�軤����/��3��̙��W<#b���ٜ�	=3�0N$fO5�kK�|��P �4m�����i�� /}垘*]:��ㅗc�s]�
Â]����Q.	�f����HK���~L���-}�7�nH���_?6�㼌th�mT6���j�H��_?�����;��>o\S�[W�b�F��=�ˣQk���hb��hԡ�C�`G� `��_?���n]kȺ�D��;j�+��x��ԉ�K��r0����6W��z^�륦k�<=�n��~����������״��A��������"��W��{oW�_�3���N��hǈ�3gf��ٵ�`��޸Vo?�+������S���#�{�o��b!�5Uj��%=���k���*������I��
��l۷o��X,�jPzz�HFFFA�������1����n 9�ׯGn�|T?`�}ӵ:;�S�a1xx�Z5��ӵO���P�ק�O�j�>'���}�����7]�W?�X�/��$JMY�~��;��f�꺽o��_��l���u�Z=��u��Ks�tq����>�=��>�{n�TinV��nS}M������ڕ�.-TEQ��33��ժ���#�~^�޻I����-U�s>�=C���r0��ݖ����{'㪜�=�ԵEya���F�/�^V��3�uin�vݺV�k��۔�f׈�#�קue+t뵫����ڻs���s׆�{��ׯ/���G�W[�����>���<U�j׭kuནQ��a��H��?��:���Gkt�z �L<��Q����c�o�lІ�Fx�+��<B���:0k�ቾKz�翉�o�?���~�E~k�Jb��tOD5N~��g�[�f��Q��Wն�Ks���e������z=��=�]�.������R}MUܣ�������k�J�|T:��U��ը�jK��Q�o�>�/,WF�~	 @8�=��}ݳ(�h��H�+�9�;�z��Ԟ�V�+[���_ZU�btRl�fk��̜j�oP#좩�:�ξ~տ�ꢙh�4Li��x����%�k��:�I
{~���|X��a�%�<�_�Չ�~}m���Hm��REa��>����5e%:��v�}ӵ1]����O��;�j2����nԺ���gS�Go\���ᾘ]g_����1�~����L��ghT�>���rm��ڶQEyq<�קW;>�ۧ{U��PuiaT���������z��.�^��FO�:uqHwT�Ϩ����麇����;��y�1W���?����~,��-U����Θ2��{'����bj�/˾}��V�T5 ;;�l~~~l�u�<��N�R� &�̽���*SS�JjY�x�+MM����bL�,9#.����[I������g�rS�{�9�	�j��%m�6���;�~���Ж�r�++�-�W���y���:���^C�_EQ�*
��N�]ZS8�SQ��'�U}M՜"1�t����̙��-U�:��v�e�����W���[,��0B�<B�x��a;Z�=��_?jHI��l�Z�}_�'�}�b	,�M�g�ߊV��SϿ~,��Έ>z��o��C|$����3>v�'T���'�YXغ�Z��dF(
��x�xlFp�պ���|?�B)  \Ů��z��]��>������h��I�t�C�����z����W�-���
sD��(O��G��{�^:ܡ��ް�N��V��{o���^~�d�]8��> S�e�1��oI��� A��a�c����k�D�%�u�����1��U����J�7_רS�S
������v��ۧ�E=ʹ�0�J���1������^��{5��,d׭kC���	}󧇴��
U�{ȩg~�֢�����+[��L�N�]ҁ��3F�������P�%�P\�#�tך?�������望�R�����ŢQϤʬ�����������d��D�����=8��!��]�᪢0O��)?ӡue%q�6�f���L��<pgB�v:������#ij{�[V�PEa��T�6$��R�>V�uh'�.i�C��X����5}���=���?���z��	�0�/$��;!��`���4����nB��Z���2?}l�IW_��5.�<�H�J�sT�]���옟c�Xd�X�i��б��9���co{2�軤��^5<�m�*��pF�����vEy�(��at"%3�IS�58�rv�x�u"u*��f/��H����v�?��g��7�r��ict��H֬r���d�Ŀ����gҫ4�'�j�ߍ����?�G��0��A��x=��H�O�����jo|(�s;�]T]�+j}�A�U�QS�5���
2jo|HY�k~E]����}���˞�#) �,�H�W�#�u~�1�R%Q�.�^��v��FB���W�����bڠ|1y���)A��SL��(O��{�*
��o��>�k�����:�w)l��p�G5��U�r�������{����g���{���W,�=c���@@���# O�P��b�U@u��'�-�: 0������oPS�fu����S=3^o����,�W�Oތ9Ѕ��9tV�.�QFf��)�)�[|ۦՋI0�xl�)<���pGB�q�ݓ:��o�>2r;�X=���{Be���[j���Pn�Z��¼�7�Gb�^���7���?c�����ڦIϰ���~`O�UzF�����R�q���X���5�c��O���O�z�Ԝ��7�q��?���"�=[�O;�W���u�����KW���-�/<��EO�-ȵ�,�@�EJȲ3B �Hǹ�*���f~��Ӱ�35J�s���7�����k�[7��z��O���h�!m�Xm��3%I%�*��9tV}���▘��L\Y�d:�wI[^80���b��ׯݯ���}��}4{m�b�!���t�����Ӫ��im�*׉�KZW�bN@���\{tL�n]Z���]j�y����e�k�w�~߫�փ���K��&<����I��ǆ���#�4��{2d:����g���뫵c}�Z�ר�'o��~��j�'�%C ���,����j������%5�>���b�6�u `2-G;UW�F;�W�y�65��MՖ���~��F����yNN���^5�xኛ�;ߩ�K��h�u�<ˬ���w�Q���3��YО׏�dDg��Ѯ�U_S�=ܹ�G�9%5o_�������ۣ=ܩ�����-e+B����:�}�o����GN�jW��9Ӳ��{�Zo�
�W����5��jxxX��.�ᰫxE���	oC0�u���h�%�[7�q�F5l���x�`�t�����n'�k9 ������l��F_x�EO�mͳ[�,ғF�S"��)�\æ�?���͡���fW|�Z]�=���ߑ=-]EJw��n��bY>�)����ۧ{��;ݨ�����K��gm�����s�}G�����j=b������E0:���A�^~�d���=��yL��~x�ywG���،-&��	�{n�F\�P��ٕ�?|����Ј�3c����B�XW�B������p�{|�����*=q% �t�#������d�    IDATu�Z=���q{��/��F����v�QU>���!g�k>?ӡ�wԆ��{��A�=����O]��������Lӛ�Vk�Ƶ:r�wƿ/����S�?]o���3U�����\Ymv�9/�\��UPP���jY,���,;�W��zMh}�l͇ޟ�~�?�Pæ��3[��T�Ԛ����>�:��.�)c�V_|j�)5�|co�U��w�&��	�<jz�jy�>�>����o����%��b���Z��z䛼�1���̑�jU 0w���D�%��{U�n]�g�ݔ���>:������,#.���~L�wLMI��Ji�s�'��[�jM��W��Kou��;qy�tO��G�{B�5��XÕ����w�N��N�vb������{u�T��U�umQ��T�Y����_dL/��j�F\�}t&��	�軤k��gs�jm��SI�s���ܢue+f��RU�-/P���Ϩ$���\�ۯ�wԆ�o����ޫV+?ӡ]���V� �1����{�O�5��j{�Ka�W޲z�v��S-�`�
K箅��[������wy�Z���Ӧ���z���{~�8I�����ڱ�zN�kj;��G��23���w��uz�᫟��~�5�[{��~k{��.��� ��h=~*���k`DMmG�ކ��J]�N�I��^�vISB�=�_O����7̎��=���;�[�s�v�?���t���=�_{^?��~��?~C����]Љ�Kz����tʗ��`��/�����go71=��>o�u|��V�	��k�TQ�7��#��ծ0[\l�Z�-aF�wm\��53�`�e���0O�gmi����ue+tǬ���j]ي9[`��^�k>�aij�qKUy(�Mn�鰇�|^v������E8�7�5���]�=�Iψ�3.j�K�50r�"&�~"Ia��I
��;�ھ�B��������}��k������� ��*��UwcE����	M��e������}���'C0�m��ӄN�
�GZ�T���k�+o�|�e��#w��)Q/�Ow���=�I���1m����m�茜�ۇ��u8�����>����u|�J��3��{/���+����<a��=�Ԉ;�}f�]��.�uI���z��M�}��՞׏���j����[uy삡�-�t� ӡ��]�Ѱˣ����V�B`����eFH#�G2]���>�ᗿ!�{0� L��������Tæ�P��. ��Z��e~}�{R�%��ͻ&imX��>}nj-�+o���JwTMM�="���Q�軤{/��ӽ�v4.Z�~���#�u��aG�"�tO�����a�%�u�IZ��T������-/���u�	��[%L}���g��qy�ďߘq<�����;Bk�z�FC�ئ�������{d��C#d�}����ȭ��}8r�W�=���33�����I�軤�_?�-U塯���P��S��r�x�==��7B#fӧ�N�{�k�v�릿�g~�������N=�ũ_���/���J��^�k1���U$�?���)+w��3c�w*��ڎ��z��nP��݆O�����y�.Co��~�5�/�k�B �PS�fՖ������t��M5j�����%�~�?��m��Hekn��s�9��V��V�#[nט|^��F�~���p%�}��� ו���Iq��3�O��m�EX*�jN�]҉�K3ʾ�*�_���<:����S��{�vzi[�i�{�\hs�`_x���:τ=���^U��8�����K�;TQ�7�ks�+o��׏�9^��U�+[!I3B���9>��h��������R�=�{n��\)|�'�.����{|�s��~�O����zo�{ZJ�N��is���3���SZUPF����;��L���݄}���B�4��)���O��f셧Z�a��^S�����:B �L�7�]#�@��YW�&T9,�i9Z]�Qc�^��=!ɮ@�+�-���IҤU�u�O�ե�C������42�*#.Oد���wΝ����FL�;>�ߍh�'��.��ْ����K��>�Ν�@��(�`�q��ר��t��\Fp�ѷ���z�ڱ�Z�[7�ն�<���@��ŧ�O�m�X�����5u `"�������4�o�w=B2X,6��W���MZ��Z�y9r��]y�*i�my  fc��U~�t�����+��5֫��Sr|����l�E���;��`�Y	�׆G��x�Oޜ*f���@@?OŴ��F_x�%��)�: 0����?�@��Ȝ�d���Q��g�TKs�++�L9y�dO�Qzf�` H���1]g�ٵb�M��s]�kt�3y'���M\��i�[Ԗ����9�k�[7���!U�ݣ.�a�'��ymyiT�	�o��}�D{�/�$�nm��F6[pyp��|�E�b��]�:#�$t/�ͦ�K��
 �Q^����^���Y�Z]�^�44����S�P_��}v��gj}�����WN_'���������F��9uk�f�Z�-i~kTSu ��4��w���C�G�bY4��e�Q8s���>Y'G��d���2r�W^�_���r����'$���� �����ʟ��V����r��S�K���l�Z��R��oC��?Sæ�9A���)�~�ID�.gk��k����y�uF$���/6���>Ց��G�)�B� 蛿����v  ���Pqh��O�d���ҭ�Ϻ�d�ov�+���ۡ��٣���W��Ψ�y-��Nijf��A��'P���J���e���N�   ��o�98��')i�Y����T�a�@@B  @d�wnU�j9ک��|Ֆ�������8w1��A��P�  ,k�?yS��^h�W�7�*�P��Ў�Ւ����k��Eiܻ��_F;zH�  �Gp�dI���"�R� �l�:  "P����?}]���uu}���T燞o�nij�)x?D�����H]æ����Xܲ�Muf���uQ���f  ��L_s5}J��a�G]#j�߬���<�n �A�  ��~�g��f�~�G���
���T7�T�O��q�F�%*�Q�d�X�=$� p�奪-/���~Iu�kTY�0�`�z KK�*),���t�4  �*��r��O���Eu�����R5l�YpS\�K��g|<}ۂ��fǹ�Qm���P����������!� �G��5顏�'s4�cW��snN K9ʊ�A�F=�*��:q��y$��%Ip=]p���������M5j޹M�z��vD�;��F�Z��RÏ~1�܆M5��;�]T��筴���y�R�^k9�*�_W�F��?8����FT����q�5l�	�D�<j~�9�g���HS!)�`��H�9�ػc쟟jMu[$��6D}M� 0��֤���B[s��W�y��*�,����Ue��(-;��X,Y,}�y4t�du��e���r;�WOU�tyB��Z?�DM��U����d:���}3�Nנ3���6��-/Uˣ��dD����T�,�t��~��n����v��ᦢ6n�0��'o2�`Q���E�����: �~߄��㲧�H
�/�2����5��f��$I�w�*v���T���h���Kp���G���G���Q������7�	{�VY����|��TS��<�,�W��m��^z��p;=��<jj;���ҩ X�F�;��� ��X,z����JϋOu���O�m�(����R  ���:����х�?�u��ώԨě�uA뇟�x-P")���v$t~pM^A�C��6J�褩i�;~�3u$Zjp��� ����BO�ӧ[����f�ێs��?M�l��ϓ�  &��%�xro��bm��RB �X{�C����io|hΈMp�g�f�M��n��?}=��*�M���;rUZ�N�׮Sz����a���N��|m��=�(S��S��s��pU�n�}��|o���.OJ�,�{��
gӿނ���h���a��8F ���b�]9�ػ#U�ϳ[�b��u ��Ֆ��Yw�~�G͇ޟ�*����\���q�b�HF�r
oP~�-�)�VNA���t��*\q��ӭ��i���,���٦����p#n�Ey��F����:%��g��CA�#�j���f�����*kKַ�&}���o��a����z���"Q��~���`�kܺaF�hj;Z�4�XGA�#4:��r��׬Յ�:{����UPT�tG��v�,KB��l�������
����N�,9��^K������_v/xn��{�0��o�Y[���:���p2������V|S?��E��'o��TO�����$��~s���TY����#	�XlZY^��kV)?7Sc����Z�η��(]�� ,N���٬�zroA�������v��=�i�A���	̷n���E5�QS�f5�ܦ�㧴c}uhzf���W�f��y갼^��m��iF�R��T�Y�[7�
�DZ�$x�|�۫�v5��>:7}�n��,�G �.����p��Ou$�9�ػ�귶��$F� `Q���-/U��H��ܤzz������v�,�����^�ˋ{�H���¯��n���lAܫ���t��Ia�x�����)������0�E��~k{���k4��O�-��Ƌ�6YfD��u �ht}��9�/���xhZ�BO�����{I	
rd�PY�M���I�:/$�ىڛ�T�UGނ{�Iх���B�nm0�|����)\x�Jiz���BdS�fISm&�0��o���=�b{�7���{�ܧ�6�٭�E	�P �\���5������a"�k��~�&''599)[Z����,�P�z�vh�3.Ir�����}Ѕ�?�;�pQ�T��7]��eO/RM�N�mܺA�;���Xmy�Zp�)��+f7jܺA-��q��r�30[p�{��`�kz�Ii $�Ţ���{���ܧ�6D�������ܧ�ט�����~�t���cM ,ӫ_�X_ڬy�=���@װ�&�~]������5u���rTV�gs��|�	Ym��y'd���3��j�Hz�����t�i=~J�WBَ���/�r�S�5�o}�k>�~�Ѻa�G�o�*�����3^�0F0c1���G�Pˣ���8_�;���q��� `f���zW�]�O���@@����uM?���Z,�JTg�h����}�: X��S�ZP-�ާ��aGꂁ@���9����u����b�)7�B����h��#��s�5��Ž���Q�h��CV�`J��z_]�N5l�	��u��Z+9��p�u���h���צ���8wQ�����nPæ�ｩ�Z?�$��1 `&��Xt�d�;�1��$}˳�۷��j�J������>���o�$�\�g:9�Ju3�����Z��z���4��}5���Rmyi�}��nPS�fu�����9��>���F�mGB#s�jԼs�T��W"j��}�Jݔ�ٌc���O٫bzO�M�����^������ׄ{0�z�d�������  �+���"�|���u���`�����T��Ֆ��=Zc�Xd�Z����U��5�/�I�E7�jK��M  `&�_�"���7����6ը�T�Z�����2�n�������oPæ�?u�i�N_��kg;?�urT�Mv�-����z���eM_)Gza�kpBҙ�� �rE��E�k`$�^���?W��ݡ���~v�װ�35%�J�pS7���/Å�?�  @��Kk�R�5u   �ǚ:    01B    ��    L�P    &f/))Y��������8��=K_q�D�   ,Q��   ���    ��u    `b�:    01B    ��    L�P    &f�t����1U���^��>UϏDFFFaFff��?�����⾧;@�N�7�M    ���/�גnJuC��>���������z�����O�    0\    &fOu ,]��"��ޛ�f   ,i�: 	㷧�U�2��   XҘ~	    &F�    #�   ����   ��T��@C�o3�*=_�P�j��G�   `g?PqW����Oߑt�a���    ��q�u}��[
�.���wT8h�h#�   @�4nݠ�m��n)� ���   @�d:����*��P���Q]�]���P    �wn��e��ڎDu�RtA�;
�    H����j?��5e�-�@T��;�H�S�9�Q_�H]��Ҿ��6    fm������d����:B]n���Wz/|��v    �lL��P���5����:9�Nus    \�V��U���7n�G�'���>5�E����f����T��^��qѰ��F������댮R   ����1�S+W(=}n����ٳ�
������46��ʕE�?�T�~��ϝ�P   `	����a��:k���w���+Q��ΟTaav�����$���    ,~������y���|��~6湉t�R    ���   �T?�E����0R    &�H   �%��%τwƱ4�_��i�}���<�3�kKK�s%B   �%⓮:qp�q�զ��I�	X�t}����<ע�Ң�<s�s�    H ��:I��}�8,�w2��1?�2��zn@}���O    �����#8�'����3#�>���:    01B    ��    L�P   `Q�_q}���4~�M#��b��P   `Q*Z���nKu3�o����wk"=+��	u    ����t�   �"�T���N"�   0���
t�   �I,�`gd��$�!w   �$*Z-�6�\:�����ut�   ���^T�k$�͈Y�ؐ&�u    �������+�͈K��H��ʨc�XS   ��B�����r/B   �Eo)� ���   ���]���P   `�Zʁ.(�`G�   �(��~��]P��({l �k	u    ���T7!��Ƈc��P    &�>u    L�s7��]��d��o�n�:O�׻|j���F�   `j��4�tj����ύ8�=:{�W���S���u    � �ΟVaQ����!��w���+1��R��?!�   X"���;/��?��?��f�
�    ���    ��u    `b��   �d�����8�f�+==mI>W"�   X">麠���Zm*+-������熞�л   @�Y�7XI���S��ay��K⹳1R   ��>>}>��|RO�x�l��   ��1R    a��7�aS�
2�Q뇟���H����0R    !�wnS�����sU���ƭԼs[�[��0R   �p�5l�Q��Sj��/B�ZP�j��vD�.ς��_q�r����ܔ�[m)\ӵ��   0\ݍ���?	vy�z�Ԍ�2T�Z]�ݖ�."~�M'o�[�Y1]O�   �4]�Ψ�_��.�@'�    ,rK5��$B    Xj�Ψ@'Q(   @U�i����;.I�w/X<e�h���T��;	ik��$B   �j�����"THe>�`Wr��K���m0,�I�:    	�q��5���h�V~�Gu_���G�   `���5�1��g?Pq���M���.y���[}�!��P
    SX
�.���p�א{1R    a
2j�T��?Q��H�X㶍��^�a�G-G;���n)����/�]Y';B   ���-/U��� ӡ�Ag(Ե>��j�KC��U�QSQ޼k�b�2"�1�   @B�<z�$����?�$5nݠ��R��T������W�q��mTA�c�=�r�������b�    n��jU�����|����su7VH�������P���4���z?Z�.���w�=6ӵ�:    �N�l9�:V��P]�u����))4�W��1��c�Ih��5>�u�:    Iz�zRܒ��B)    7|�-I�,�m*�c}��?�������nX��6W�f�?޸�u�<�w?�4�g,���F�   `��h\��jz�*�th��ju������.�<@s:�re����F����=۫@�؉��z�l�:    ��8wQ-G;հ�&4'MU�j޹Mu�kTY��+CL    IDAT��������u���
��e��Q��[~�_�Y}����	�   @B4��Mu�h��j�<j=~*T8%8B7�����3�^����;/��?��?��FI�s��    $L���n*>���G�P��S)h��B�K    	S��PS�f�U���Z��j޹-��#u    ���T-�ާ��|Is�T競�T;�Wk�~皺勑:    	Ѽs�*��`��ޜ�+����vD�5��f�3�]�pi|Ɵ��IC��+1R    �ר����EP�����5nݠ��5qmL�I���88��jSYi������zNB�   `Y���B�B�.,��&Z�V�����wqX^��#g�z�l��   H����50�3>>}>��|ROo\�Y,ϝ��:    ���`���ω$ b.B    ����X_}�s��P�26�:    ��8wQ��O�q�5n�0�y���O��U$e9cM   ��h�ɛ�,�WS�f5l�Qǹ��tJ�*��T[^���|u�����6����m�ڏ~%�ߗ�'�Ǒ�K�T�t���,Y���[g��P��   �IA�C��6j�-7�Y_�50��?Q��i��	{}���%�<�l���ޘ�'�E�P   �'82'M�H��-�`o���~	    I:�]���Dz�N�|��vF:�P    
2Qo&��q���0�Z�3*�I�:    	Pwc�Z�/�k~��?5��K%��$B   ��8wQ͇ޏ���	����bmZ��Z�r>J��R    ,Fl>    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01{� s����5=�RZz��2?�_#���T�   0�q�8�У���T7e^�/_V mT"�  `	b�%�666����T7#�˗/���?��    ��:bllL�������������@��   $��SZZZ��2::��&    	G�ò�ZT�e�l�,G�N��   +B���4�ʍ��YRR�����a�   bE�    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &fOu��
3��ސ���C���ci�����|�c��n  �]y��+�R݌��,�zzc�k��
=���X
c�����f  `W��T7!*�:,�>cC���   bŚ:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L̞� �P�f�Ck��_Ia���/v?    V�:,�t}�q�%9��   ă�    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L̞� ���Kg\~����v/    �:,�~}�g¸�\2�^   @�~	    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���S�  rm�Zlܗ{aN��߳#��   ��n�������F\~C��?i��%�n�=����\B   B�2qflB����o֐O��   @�XS    &F�    #�   ���    ��u    `bT��i�|>��n��~�l6eff�b���Y   @R�`J>�O���
�$��+�׫��\�   ��_�nw(��|>MLL��E   @j�`J~�?��   �RE��)�l���   K�����)�u�oZZ����S�"    5(�S�X,������D��%�   ���e�X�p8":�������۸�|θ{   q`�%    �#u0����R݌�ݮ���T7   H(B1>>����T7c�ϧ���T7   H�_"n�5�I���S�    a�C\&���-(UAIy��2��_�Y��n   ��:�er�u����W5��    	��K    01B    ��    L�5u �����A����n  �p\��&D�P ��seU��  ����K    01B    ��    L�P    &F�    #�   ���    ��u    `bl> �jJ��o�ָ�:����g:�t/p%¡? X~u R*7=M5��r��c��e�m)l�yџ  ,?L�    #�   ��1�@T�\�*�՘˘�YΡl��������\.��*��D���ONhrx@���2�{%B�k\�?9��˗��Ŏ4��o[���CǼ^�F�n����}�I�Kc�C�>�x��  ư���r��VZ�����+*��\Y�7�\s��ۍz<�(���u�~-��-��<E7����ؤ���T7e�  a)��:��~(�m����T>0���n���oVVV�$���L�C.�K����$��ŋq?o��d�gFF�._��,� ��lY����<���'�===��'�a��7���v�r�-��?�3�p�*//Waa�$͘&8��������&&&��ե���9sF��c
&�%�,������ٳg�D ��-�PW\\����<��?�?�KA�$##Cw�}�n��v�|��r8��H�|>���kddD:y�~�����O?���"�'  0��`�C�xV�������l|��SFA���Mx������!MK�XȪU����k�ƍ��Ϗ;x,dhhH###�����~�;���Gt]���	  �Pg����r��p�je���z�r�\���]�����٣_�V2��4��U�V�G��͛����@ ��VNq�\�������~��_GF�Db��G}T_��Sڟǎ����z� ��Y�.Uk���Ҕ��-#u���x4::�����s��r:�S%�P��&�dggk���)	s��\.}��gr:�:x�;����
"�'  H�e�R���D���JKKKe3�˥��A�^�z��������'�۽dB]��n�����׾�5egg'tZ`��N�z{{500����/X$�A$��|�ǔ��C ��-�!���C���EVV�#u&�~�����y�������D��$�.q" ���z��'��C�f��t4)�á�������v[(��SPP ����ߖj�4�����	  �[�i�P�x,�Pi ������|G��r�|>_[�ժ��Y,]{�*++����Þ�� B�  H�%�6u��ru����K�>������h�|������)�á�7�>�����"�'� �d�,#��E@�mۦ��~ZYYY�	 A999���T~~��y�egg�=���R��O���b~��'F�'  �:B��E@�|�ISoϑ���믿^iii	"��\;  ��	���������T61p���ʕ+<���������Ą�_.� 2���ҙ3g499�={�h||<�y�Vq�?��O  9B]�|>edd��΄&''5>>����ϛ�������7U��4��]�V��������$�.�Ad``@���w�=/� BN����VSSӼ��  H���b Q�$���g�UVVV[����*++Sqq�{�y�N�����9՟��'  ��X�2�� z��'URRb�"�*,,T^^�jjj�iӦy�+..�Ĩs�{џS�YXXhH ��� �q�}���n[������L��k׮y}a���5�\#)��	  f"�����Z?�pؽǖ�ͦ��2����'�H�3�[�Y�&��	  �"�����򗿬���T7%irrrTRR���r�[���{/�����LX ��u B6nܨ��k�O��k����Z��G,�Oc�  �G�K �Ͷ$�X,Kv'�e-##C;w���MuS��f����D^�W�a�=�Oc�  ̏]��b�hrrrɭ��Z��X,���,��V�|>ߒ�����jݺu���HuSR���D������ׯ���G۟  `~��
Kr��|��n�+==]�E�@@~�?�-C��v��o߾,G����K###ڴi��=��Oc�  ,��0�����˗5>>.��#��*�����5�\�[n�e��"��n�q�q݇��bT ���>�/�$��jbq����+�����)������<]w�u*--��>����  ,�P��
r��r�\��wX\���USS�$�
�"??_N�S_��c����)��  W�O�H
��/�˥��IF����UWWS�押�<�|>�_�>���ϙ��O  pu�:$���._����ȝw޹��~Mg�ٔ���իW+;;;���ϙ��O  pu�:$] ��c:fj��v]{��Y����v��nݺ���?�������X��	  "CiB�������f3������:+oKQk"������J���Ѳ��u��]��Q_G�k ���R�gI;�ͦ�˃�nF�


�f͚e�A�|rrr$I7�pCT�џ��ڟ   2�:��R	vf�j�*
z�#--M���Q]C�/��  �aA�ǣ@ @�$#����p(///�k����ҟ   2�:,���<�iq�+--M>�/�>�?�K ��갨�\.��K"*5�/==]n�;�u`���b�O  ��aQ	r��
)�����jrrRn�{��&''�!   )E�â������NA   ,Z��~�=`�w���Y��X��
��b��D��P�EirrRiii���LuS   ����7�����w���?��X��m$�ٚF��,v%j��P*vQG�W�΋�焯jܽ�(�!,��=lv��E�[���L���oþp�C�2��]j_%G�nD'e,%��&��-r�^P3�(��ΐ�~���4���cZ���{� l&r���Ƃ�~�踽�b�
���Cz��I�;�Y�2�eɿza,\�/�ŗ� �@ۙq� �~��;&udZ�t��:"�K�����n�0��,�?�����x��/����u2��u�_���Ů����,��?h{��X��v���Q-�`�K2�Z:��j����Қ��Y}��E���Ç��Ԅ۷o��1���ʙ�z������.ڛ�����8��gB�Nf�g_�_�y�,c:-Jn�:�ű���Q_�	Hh�� S�d25q���ں�k��L�ϬVVV��imll�b��4G���ʙ�zu�DU�?w�/!��2z �^'s{��S�1�����WǦ�����PZ��Z$v\~I��N����Oj"i6B*�*yo'糰r�^��_�k�o����Bu���y�4I��dV���+3������X��EI�:6�rn�m�İ t��<L�X<G*���e�Ւ�d����d2Y��8�;+w>�ٕ����P��ש��@"��<�H��WǦ���Z �U�s�#e2�ZY�Y���8��鬭e�A��Ζ�8���ʝO""�j� ySǢՎ�r~,$�}<���2�,��èK�D�h�Is���U�۷��~I��|���$""�&YƵ��c!��/�%���x�A����_��IH���U������|����<�̧����=""��TF�:��cqY�|�<�wT�GI?��կx`�L&���|��Ge=�����|�t>��v� pr�β��Q�e�̈e���/�˩�1�#jp������e�iii	{��){�W<�|�t>����A���c�,��~I5A�$��P�VWW1==�g�y�t���.�H������/�z<�s�T4�fao���œ눛��<=��ن�_���{��|�'��}������� G��� 89��cO�  x.mm`:}ng\���h���'�կ{���:^ṕ�7�r��u���W�cj�����ف��_B|-�_\�������9������?r���7��Kptv�s�-�#s[����q�?�v�^Ͽ��焫�K�Z��M&n�<u�#��R��ւ$��K�/-J�=�8Z�c��QM��V��������6|uiccKKK���X]]-�y8�YXYY���|E�Y�o��#��@;:;��4k%�{�����\���y\җ��w����7�:}����������7��<�^��$wv��:  <{��mq\�]����9z��7կ��=�n�w���I�u�f�/>���|/����aDc	�[���-�,N�xsW��v�d���x����W����z�����\���Ww�#��� w�͒?�*�ukFF���K�:6�~�b��s���j�,�쀩�{��arr�����/���}��������|fi5��8:;��߮��;ث~R�5����]�(����w5�I�_K!89O�S�R�G���l�;��0p�&����V) `j~!{��G��;؋xr���G�_wtv�7�Z���:�[��(�����$��������]=��ȅ�#��QJy��d���ϏB[ө�x_[MZKQ��֊,c��w��D�I!�N�ʕ+��d2<x� ���wiT��jm��ZΧ�n�Fpr���7@T��k)����-����!����a���M���ݥ���~���A|-��{GIDɼr+j����|�X��7���U�>'³w�u�f[Y]{Ky�+�'gv\�,-ͭL�F��[+�(��l�JM4�� ࣏>���߰��!�"���I���裏��{�5l���|U�����^�g� �ހۛmE���g�l��M�/l�u;{05��pdnK��݅����b::;�Pc�9y����jUMY������E�Z����lC��mDc���BJ}�k]iε��M[5���TSA�:��������7�7�,��`qq�dR�$d}}?��Op��Q�g��_@pr���C!O�n��$ `oi*�9ów�*���)7��X��.�#sp;{v�KUh�f~����S���yy��L� ��f)	X�����u�N��o���5��K�b����Nv��A���BU��_����������uki5m�嗒(�E��u��3�������D"����w��d2��S5��9�����D���|j;�;��4!pr ��H�^%1+�r�U��H���7���F)��I�J���CM�����Dpr�`���F)J�{����եQi#���MG89�Vn�#sN��7<��q
een2�u[��۟K����L��N<u��%��zݴ]c����ӨKت-�N�ҥKX\\l�����
���055���/Χ�{颱��u��=�})���%�?+�U��(��q{�S/��ei��d�ꏲG�X�����rM�1�����-I���N醩�2��Z*۔�ن�<?�Gm���K������J[.�<�xr]�v�sn.��V�s�����J}�Gc	��b�[k�V�tR"Qݥ\�J�.���X,����A,3z8������O?��������|�'p�fիc��&8:;ؐ��'gԆ��	僃��������V�$N�����Z
���E��q�G�mk;O�S*j�+׷��
�:���E��|�':}b[�47�*�� ����RI+t]9˗�zݴ�:�	�R�0�p8���Y�����O>1z8��x<�믿��9j
�'Q��_��M�N�@���-gw���|M15��=�+����=Ww���J+��BG�7ԏ�t������a�Ȍ|���N����Y����t)	���+{v�G�($=}�]�J}����.1����䌚�z����n[Z��^�6�ba��AJ�2�#�mdY�ݻw��3�`qqKKKFIs.�}}}�Z��/̝�D"Q��jΧs�؞(�P���\  BIDAT�)���\z+[�x�Y�#_82���;7;��t�������#�N
5J�M�	��	��4��f*JI�vJL�%������<�_��]R�YS:izLh:�����;>�����^���|C�p9��1�끫7�<����׭�R���.��:u��!��j�j�8�r� @Ū6�H��X[[C[[[��666 I��կ���s����E��{wnWl�o����G^��ֆ��&���u��9���Kx����o�vyy�}�[XO����p>����
�����+�������������/!�+��b�`o���+�!Kd�[��|�'���qQm�����Q���P��w��_��V���,����hH���hii�7��M������0zH{�'��/����ʾ�\���ػw/�S'�f[v�[K���t�;jz����� "�mб��g��X�� �U��>��/�����X���Ckk+�}�Y�ٳ���T�'����Eww7~�ӟ��+�q>kH|-���f4��c������Sy%"jD�\z"�#o�`��L�	�9ܻw���>[�&3% �������B��7��>rP�6:5��{#b��߷��;RǢF���̸W J>��I���j��ޝ�����~�ݻ�������n��	s�\�����'�|�4	Ƚ{����Y�����i��ԛ��R��WΦS����g�N����v|���|�'tI���ID�a���JkP���q� ��rʤ�L�V*u+++��ں����yҠ������hjj������֭[�����\���nA�$�A���E,þ}�jv>�|���z��&�`Z����o����y�Spr��j�o �'������59H������}�`��{N�@��'{.���\zK�$ˈ�Dd.����[�n��T� &udb{��a�Z__������o���|��)��v��N����x���ҎVVV�L&100��,Q4�@<���g��r�O�WTEs;{�9�=�|�\1�ȱl��Ko!��B��	�G����F\�]�N�;Ҽپ}�Ͻ��V|��1�ȜD���s���cSՌ���G F�}<�:2-A I��àH��h4�'�|_��W��_��Tg���v�����~�3�/�$	w���|�(p��p���D4�P�y�7����BprF��g��?r��.�Ԁ��5t���ߏ����lI�k1&�� tX3b��n\�W#f˹q�(��J��I���je��ܽ{�(��v�Ν;����L&������׿�u|����/~a�X���ԇ����%s�{����;�״>>����%�k���*$v-��]VI���R���Licc��q7J�LX__/z]:���b�Ҩ�I�ڵ��bdd�H���UMF����tbqq����*��,���	�P6��;d\�����X����<G#��ڒ$���_K!�,��B��ē�L,��4�$v�s�^��b�;;�%1XiB0�#E���D#Hg2�WCWWW��'�����'�O>�sss�{��f1r555�駟�7��M<��Sx�����Q�8kkk��Tr>wo7�[ng����-�=}N ����b��U�D3t�6|��>�ݯ��H#������`/<}�-�5���ݲ�3x긚P&n����|ϥׁ�F�$"��Y%1�v����~XVW����7�����.�:2Q��5��$�i�^]�������������a�Z��"�U��455��p����~�iX,ܸq�n��h����q�=t�f�Z�900���fD"ܽ{�n�s��Gf�g�K�#��������	'g*��4D�S*e�/4ѽy��|C����9�Mb�Rj7N��1 ���.���b�<�݈�DT�C���3=A�W�|mgƽ� ���FC �F��2:t�m�Z�=�=A�N�M��/�� �J�����u��˶�6����������9Ċ������!<xP�f4� �w~�w��҂��%ܽ{���H&�XZZ����n��n��'�@WWzzz��ގ��ܾ}��_^^�.�����c_)x�Q���c��/����l���`�����a��=p���l%+pr���o��{�Ww���SO�f��ܫ&�J��WA�:<u��v�A�>'��?�������VFDD��2�ɐ���v���6:��k�xA�i��)X�#S1CB��<�;�{�H$tODdY����YEtuu���v� ��������b�ǿ������}�>��3]ǘ/�L"��m��!]$���OeNͧ�b���>|�>��ABWL��M�:GgGv��?e_�w��f�nU2{K��6�5�#sۖ*�A��Dc��؛mjsV	��A� �+~,��xM�� E%���D���nA@ �:.&ud
� `mm��a4����o�z26����ê!������qUc���C,..b5��M@�������AI���:�sS��Y	-����=�F82�m��lC���o���t@�b�v���Ec	u�`82��tD�`˾�z`D���jY�F>�c���<"2� �9A�s�q�77��*��dRG�cBg�ŧ~�O����֍5H��t&S�18���G��e?���~��}�6���#����@ =��.y���S��Ep>���n�[�89 [U�7���_�xo]n<GgGիb�+�|�yO߲����D��0����߈ʕ��e����VM�}?
��C"z$&ud�zI�������o=��-xʰ���_��aߖ�#��8���(V�W��많j�4��M�g!�X�����;5���bGg���������*B�x7��^Q�2K��7���@��k�臈�:2� �$���ՊL&����F����ެ��T1ng�#�Ԋc�A�z%t���-q�J��\U;���Tٿ�r�!��7�`oiR�\��S�LIGgG�^�Qg[*��Wy5�Y�L��,R��.�߉�1�.������S7�ă�3�7���s"x�8��?�M�n���FШ����\U;�����lSv刊\�X�n>����;ػm)s4�@pr�n^�"x�8<}N�g�����I���z�5��]��=��9�f���}�M������D��_|C���;7��*����	�8z�hL�j!�S4�LB��� D�c��fXͩڮ�&�LWw/Z�h��TZ���*�ĵ�x�����9���8�Z�J�����s�7< �� ³w����X��Q�2�ZO�#�\�~8Q଼hgG]$;��~�G�!�C`�Ɩ9v;{����K�#�gD!Z'�~��TϷ��"�{�������c6϶T��*�� x���:}���۾noi��ϩ���~���^�瑲�AY�`o�m���^1���`u�
�YH���F�n4�|O���A&n �S[�+7��Ύ���t(u4��c���j����_�6E��O�3{�����MGt��f\#*WFV���;eI�N�.��3�*,��=z�>�#�S:�j�;؋���}�u�x89�k�LIr<��R���7���^�c�ów�9�mń�ϩv�՛+?�����f&u�+�ł�����;GD�|�}��m#%		��<|C�e߈���[Yf���;���@��M�JN��Q�j�j��r�\,v���I�J�� �U�Bϭ����X�X�����v�Ճc��s14�.OL�4��� L�y\�������͹��_���S�!�֢���oX��k&L�Hs��$1�#"]){E
-G�7G�~#�v���P<�bdoڪ�߬q�H��L�]�]��>�z�S�u;���P�Z]Wx��w�S��$W��٥�:�+�/�SϑT~F(U�����ȏ�z�5�{ng|C���sh:���F��	&��z�;ث~ �,�MG�+66_�s3&uT1Q��(�2��4R�����r�����rtv pr����_���zc���ܛ&=؛m�A��.u9dprF�O����/�8�ju��FLGgǮޣ�R%�_���q�i����4�k)�.OTe�Bٓ:}b����t����^/��_|��
��]{�������h,ϥ��9�.�ԓ�G!��=puw��ݕ=Sts�|��[��}�m]�`�*�q^}�r[�֫F�A�$X,�AH��l�,�2$IB&���$.�� �J�����u�t��(b�?�����vS������>�]N�s`w)��6L��7�\�u���O�7<�h,���}⮴�w9 �7)1:�"prX���	RDc	]MSI빂��܎�
e?[�+�
=�*U�|��l��Ko�����<}N�g����U�yV�{T:�V��7w�`�_�QX�����2��٣V���H;��|�o�Om+Y���tz.��pd�����g;�uv�]��v�d+�U����N�����}Z��3"&��B3��ԃҡV�_֣��N�7��5?�^{��6ڛmp�oG���sh:�=Ba��g5��V&��z� �1�#"������P��ܮs�P�JwKe����U��[pr��5=.Wi6�׍��g/�S ��<e���/�Sa�� �����+��_���wt�˸�B^[:?�eRGDD5���;�޶?G��f���;؛Mb7�f�S����B|-���͓{�m�YO��3�:(���Q�J(dj~�>'��ܤ3�Q�I�R��=���O��~v�2n�Q:��/�����.O�庺T2�|$=T��?r��~� �h,��郒�j�`�[��N�S���g�s�<0Z��s�'�y��LUc���i�9�������Ҕݧ��Z��p�e�Z�k�܄`RGDD5J�\�$����W����-V��(�l7��	\�	���j�,����ϩ�M�!�@v��w�WӤ.K��YT^_4�@0�:���P?��՘�u�����S[�+���
θ�k��F�O� &uDDT������r�Զc�����vـ����-M[lG�%��^B]���+���[�##�#s������Mh�D24��x#bc�9�z��89�P?B��޻�˸�h�����J$�~Y�x���r|C�r@�w���c��!ttv`�� |��[����&s���e�o�_������j�é��TZ�m3"f���T��z\>���P�V���.O�t�q��J� &u�bRW�����(	�rV�B阨Wg7�X�l� ���%L�����|C��l��=�[��4�<@3P�*���qT�2n�)��L�t5??Q����F �22����+�eYF[[���ˤ��teo�e�gy]7j��r��;��٦&����S�SL�`����^�r��ۆ^�3.��j\-=*������?62<U��?��Ƥ���H�0.��z�J�&� �$""""�0�ƛq�lv���~IT3d�daRT���([\� ; �-�3h�DDDD��R:�I���2�ɐ���pq,^�Ұ�l�㎽�Gd� ��DDDD��R:�I�)�2�eɿza,\�cSǢ)   �vf�+��������L�LE�,��/�0���-_bt<�n�0��s�QG����O�����G_ȸ�˸��5J��3��w\����������x��AU�~�k_S�<�9u5��s�V�&���2��ɛ|ul��'*`��q�1( z<?Շ}ˋp����� �2���D�c���#�U������f��f�1��A�t�,�����u�$��x��饌�ƅ���*�r~,�rn�m��0;""""s�4����j���Ts+���ș4�)$�[�_�� d��XJBW��&���M1�#"""2-:�I��$�3���CF����2�H[$���|�WǦ���Z �U��DDDD��V	� Iݣ��E�~{�Y9?j?{�"���nH��t:���	��={�0.�2n����q�;��L�J�ؑ��2��\)-�ۭ���0�QdY�Ç)$�Ɋ�KE8�2�G���q��Fi�yf����5�:����O?�4�{��w[!^����R�k� .���3�>Al�8��A��bEKKKE�H�_�V�uW�D�q��Fi�yf����%=: `[F"�2~��85z�Ƃ2�0zT�_����ʸ�˸Տk�F�gƭ︕�+���B���c�4z T;��E��/P�e\ƭ��N�h�̸��\z&t@/�$2+H��7n/]��(�H"�ЮY,V,..buuuW�>���(�2.���m[��3��w�R��LꈪOF��!�J�:6�~�b�S���)���n?����q�v5�<3n}�ݭj$t �_U�,��G<��M"""�ZW��`RGTu�(��C>S&�DDDD5��	��������H3�N� &uDU��6_Ǔ�C"""�ZcDB0�#"""""҄	�����Z�p=�|�$����IQcRGTef��	����DDDD�;Lꈪ̔	� ��C """��X� Q�1Y�rn�%H�0zT[�v;���vumkk+�2.�(�Qm�����:�*��}g�=+��BF� ���5zT[Z[[q�ر��J����ʸ�˸�5J��3��w\3��K"���)������ڊ��8��V�'��˸�[y\�4�<3n}�5+&uD|�6:�0zmgƽ���v��_��r�2.�2n�q��h�̸��̸��� 6�L���u��vA�ŧ�!Bſ@6�@v��2.���(�6ό[�qk�:"��3ro]�U��JG�!�"�V+b��2.��X\�4�<3n}ǭL�$B��w'_��f�}g�=0Z͘T�dY�Ç�q�����q�;n-��:"	@�5#1:n�V̖s�.b�Z񈈈�H_L�&�k���j$v-��]VIs�%Q�`RGdJb�rnܥW�}g�=L興���`� jE��q��U��A�M�,��/�P������ͦ(�CG�����7��O����v�e\�58�Qm�����8?jH~Ťn���Q5�2�eɿz~,\���
���C�����
0*�c�K"<g�x����k2��r!\��汶�q�^��#���Q�cRGdb�����uX�c���k��0)*	��^'�� ��p� ٠Q�1�#�������G�f��DDDD��/w�ҽMDDDDDT�d׌�ͤ���i��@DDDDD&$`ʨ�L�J C="""""2��(��ͤ�˙LPF��������C�q-��+u5��X\��ݡ�DDDDDT�2��72>{啡��ũl�x"""""jd2pq�����1�RW����f�""""��&���L��sq,���ֶ��������Y��=��/+�v��|� ������d��$��αfR���q{���L�������|
 ,A
��=�|�����I
    IEND�B`�PK
     ���Z$7h�!  �!  /   images/e0155ecf-753f-4e63-a512-9d8bb2c3e0aa.png�PNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK
     ���Z�j�7q 7q /   images/b909fea3-6005-4c04-81af-b407c7630414.png�PNG

   IHDR  �  
   ��N(   sBIT|d�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<    IDATx���yp��]�������j��������cB`��%�I&�����c��0�28CXc&�0$�0lEB��P!�YH*�,l_�����-�����rt���<���s}��O:Zޯ*�9:G��~d����}��       �#�^�O�i:j��u�MH�z�G��5km�{?,)�4*�x�����$+���������T>����^�-I泼�%�6��%e���c�\��}����u�:���ͽY��kIʌ1�ι�1�m�ْԶֶ��KQm������M       p�>ۅw        ^�J�r&˲k�s�a�ix�%�{�G%K�T��״[*/y�cI��>�^i�{���C�W���rcL���H�i�lߑԖ�-i�Ӓ��_6�4���ι�0�������       ���       �Ca�T� �sn�3뽟����OJ�ޏH�{�+�-�G�,�tH�
���}cL����)�Ƙ5IMc̲�~1�{��[�~��vO�       �r�p       ��Z��:�����1��~~�D�)힪>콯j��NI�d��ƘT���c̖�uI�Ƙec̒��N�/Yk_���Ypd       ��f       #�Zm&˲�s�]�t�{NҴ�)������/y�G�1&7��1mc̦�I+ƘےnXk_���O���ꀣ       ^#
�       pT�չ<��L���c.y�/H���7�J�e�}4��qe�M%u���MI�Ƙ[���� x!�?�Tx       <
�       p��(�<I�o�yz�������1�}�{{���1�cc̎��1f��h��潿j���I�|b�9      �$��       �3\.�ߒ��%=�F�y�\CR�{_��s-8A�1�1�k��2��3�\3�ܒt5����$x       xr�T      �W6Z*���{���7x�/z���#�����:�IǱ����(��a� v?l� }�1VQ�X�(�$#�Q,I
�ݯ�$c��(z�'
C����Va~�<E��+M�O{-�29�}��\Y�?�o��4�$�Y*�r�+�ryy�I����S�;����,˔����4y�^��{�}z�1���[Ƙ%c�c�'�1�����5�       pTQp      p���ι/����ؽ��ι!�}��� E��(������p��p�y��zE
�`�q����;_����\i�*�w�i�*I���|�,˔���4U�fʲݯI�^K�DI��{?�o�H3����������{����:#       
w       �A\.���9�%�����?��ޏ9�=���֪T*)�c������()z�׭� {|J��J�
�i�(I�Ǟ��~�W���O����$��%�Z��;���1���?EQ����G$e��       ��;      ��"�T*�E��_b�y�����~�4���(R�\V�T�-��v���e�⇯��EV���ޫ��+�'���z��^~���������97�؇j���������+������?      ���;      ��f8���������������t���*����J����RI�rE�JY�RY�JE�rYA:.p��$Q��S����u�{X��������t��uO|��Xkcnc�I�q�����ʠ�      �kE�      ��T.�/�y�$}���)���ܸ��D3�*��*���ժ�岪���c��J��J�� 8�����t��u��t}�{����2�o�ٶ�.J�e��������z��      8b(�      ��(��s��~�{b�_A�Z��j��j��j��Z��r�S��8��$����{��Q���N���ǎ���(��߻Ƙec�U��       ��s�      ����Ev���ܨ��:�~cT�TT��֫��^����y�TtL �ޫ����N�S���v[;;m���(M�A�|b�P|��Ag      p�Qp      P�z�>��������޿�9w�{?|�Od��X�z]�z]�z]�ڐ*��ʕ�FF��#8b�<W���N��v���ζ��v�mmoo��1�[k7�1��1*�_�i��$�:      �����P      0xQ���ι?㽿⽟w���ʃ P�>����GE�Z��zm�y����������������n��no���V��t���㬵Mc�Ƙ?1��~�$��:      �㇂;      ��b<���I�j��[�sg����t*��V�jU###Q���evc�ͷ��sΩ��������7�xc̖���1�Ƙ�/I�ߖ�5�l       �6��       �4�ju6Mӯ����g�s�ι�A�z-����𰆇�544���!��C*�˃� ����N[�[���������������n�;�x��Z�7�,c�T҇� ��~�}й       �     �S�R��ɲ�/{��{�f���s�4�\��R�|��><����2;'�8��4�-�ookkkK�[[�>ϲl��>+c���6�1/Xk?$�%I��A�      0��      N�r�|.˲�"髽�or�M{��A�z%�ZM###��訆�J�a: +;;;�����榶�6������-%I2�h/��Yk��1j��Wa�z��]t.       ��;      p����~�����d�8�522��e������T:���DH�D[����ͭMmnnh��V��t���c'���1��r�׷����      @�(�      �_5��o������;�+:�ˉ�X�z]�#�����FFGU.ɸ pj}f��@�VKY�:ڧ��v��w�1l��`�$���ޠs      xr�     �c&���c��9�e�����||Й>SE���i�Og��냎 ؇n����������666�t�G��[�ڛƘ?��W���t&       �w      �h��q�ιo�޿�9w�{:�C�kll\#������j�ڠ� I������FkC���6Z-ml��$ɠ�I��1�Z�4���1�i��ߒ��      �ˣ�      !�J�K�,{���K�s��sG�)���>>���q���ktlLa: �����[����9�X�$km�Z{���~5M�?t&       �(�      ��q��������Y���h�A�ѱQ���kll\c�c��v��  �X�$�h����j���͵w���1�#Ƙ���?��h(      ����      �z�>�����{�_y�?�97��5�0�46:��d�����Rf ����Zo�k}}]k�U�Z���ލ1��m������� ��n�{w`�      �Sd�7�      ��*��������+�s��s�Ag��H�������54<,c�T 8:�,�F�����Z������ޭ�;�ګ���3��R�߿:�0      �	�]+      � Q�Yһ��_u
�QibrR�������� # �Ĳ4U��҃�z�`M����XcL�5ċ�0��n��၅      N
�      ����-����s�s�4�<�z]��)���kr����1Nf �h�^W�ֵ��=�}mmM�~ Y�1�������A��{��$      p�qw      x������y�N�ܗ9��z�Ae��H�j4�4>6��FCq*  GF���Z���ZS��z����s����Yko[k�M����>t�!      �c��;      �Y�q����o�޿5�����p9�1�����5��"
  ǎsNZ[k��\UsuU�^��sc��v�Z�o�0��n���C      �     �=q?������s��s�A�(�+������� p ?�}���V�%���f0ƤA\3��Kk�����5       pDQp     ��U�զ����$}�s�sQh��jllL������dC�Z�c  p��i������ִ�l���5eYv�/�A��z�ۇ       8"(�     �4��8�+ι�{�(�����&''555���i�OL(�Î  ^��^�ֺ�ͦ���j6W���5���c�����̲�g%�5       0 �     p��������;��K�ܼ��P���a���I5SjL6Ԙj�Z
�  7�v[kkM5��Zk6���yh��1�֮c��Z�kI���C[      2
�      8QJ���ι��{��<�/{����F�&&&43=�F���	Yk3  8�nWkͦ�kM�5W�j��?��Ƙ<�ƘZk���_?��      �!��     ��Eѻ�����\�\�0��J%MNNjrrJ�33�1\v ����z����ڪV�����~h���mk�G�1����/IJm9      P0�     �؉��M���8���sn�{h׹��SSj4�49�����a�  �H��Ssu��	�Ux7�xk��w%�T��9��      @A(�     �8(EQ����8��r���W*M6���U������a�  '������}�5����<��Ƙ$��K��,�~VR�P      O��;      ��(������9����R������jzzF�Z�0� �S���heyY�+�����^�{�;�1�֮���3i�~���      �w      qE��޿�9�f�\�0�c466������kllL�p�  �v��X�}YI��Nkm�Z�Qc�/�i�I�|)      �*�S     ���T*�y���9�uy�_�����[��wOi����쬢(:��   ���^�V�Qό�*�܁�4�xk���A�{���]      |�     p����WdY�^��W�y>~;+����g43;����˕�X  P�,˴�����eݿ_[[���Z�e��wA�l�����/      �Pp     �A��a����s�Mι?.=M6�����̌���G  p(z�������xO+��J��@�Ykk�ǌ1�����I��B      �j�     P�����~���<���?��P###�������&Ap�+  �{�V����e--���ښ����㭵���������-     ��D�      ������w9�ޖ���A�Vk�����̬��gT*�z%  �������|_������%�z{�z�Ƙ�7��H��=�e      8(�     �����Ȳ�ι�v��.c�&&'5?7�ٹy����:  ���Z��Ғ���������n��Xk?��������     �D��     ��#���۽���{�s.:�ea���i��-h~a^�r� �  �h�~_�++Z\Z���=%Ir`������O�1�g���,��2      �(�     �j�(������y���{�z������ͫ15%k�A�  8���j�ZZ�+�����.c��ີ��I��oK��2      {�     �r�Q��{��y�����Z��Z5��4?7�������Z  �Ϣ����Ғ�/-jyyEy��c������ג$�QI�Y     �c��;      ���}y���9w�{`׎J�����5?����EQtP�   �:�y��fS�K��{綺݃9p}��~�Z��R��v��z �      p�Pp     8Ū��\������<��r��Ȉ���5?����Iå)  ���{�V����E--��������+�ߵ���R��w��v�@     ���."     ��3��w��~�{ K� �d����-,�Q�Z=�=   8<;����xO��U9�dO+��ߊ��wvvVd	      �$
�      ��X���+�_���u�R����-,������ 8�5   8����������+ϳ���^*���n�Wd	      �
�      '�h��0J�s�:{�ffge�=�5   8��<�����i��=�z�ٳWv��i��_R�@�      `�(�     �,�q�A��k�����왳����1\f  �.������;�{綺�n�;�1�Z{3�_K��G%�_     ����#     ���q��<Ͽ�9w�J��z]s�:{�&��X  ��{�V����Eݾ}K�[[��0�� �c~>Mӟ���      ���;     �1��ۜsߛ��z��A���:s挆�Gb   N�V��{�����;���,|�1&��Ƙ_H���$�      �@Qp     8FJ��_�����s_윋b��ȈΜ=�s��ihh� V    j��ZZZ��;��l6�o�ɂ �� ~����N�      p (�     qQ}�����s_�+�qn����Μ=�3gΨR��   xE]v���������i����      �0�     ��r�|>�����/;�F���x���ٳ*�+E�    ��A�݃ X���fE?��t�
_      �}��     pt�a~�����<�X�pk�fffu��9��/(���W    ����ԝ�wt��mmnn>?��A��$I> �S�      �n�     ,��9�7��/���"g�I��T.��   ��e�۷nj{{�����Ƙ�N��g     �ׅ�;     � DQ�g����{�s�R���K�gΜU�R�x   `�67u��ݺyS�n����ھ���a����}���      xU�     I�RYȲ��y��sn���###:s��Ο��z�^�x   ������ښ�ܽ�;�o���:�Z��o�q��;;;˅     �ˢ�     p��(�����<�{_���;w^gϝ��  �S�9����u��--޻�,�
��=c���e�ߕ�
     �G(�     �(���{��y���>*rv�Rչs�t�����9   8�<��EݺuS����\q}tcL�G�0��^���     �$
�      E����s���|���Qi~�Ξ9�ٹ9�e   �H�Dw��ѭ[7�l6�m��
��K�����v��     N)�     �S��p�}O��o��v��Z���Y�9{Ng�aQ�  �SiggGwn�������.l�1�Ap��i��da�     N!
�      O ���x��W��W:��"gOMM���:s����    �4�MݾuSw��V�$�͵�����k���$I>Y�`     �S��;     �k�a�>��{�<_(rp}hH�_��U�Պ   �8�kiqI�n���Ң�s���`�Z�+i�~��^a�     N0
�      �"��/�� ��?�����3�p���gf�   �	%I��w��֭j6���5��A|$����v�����      'w     ��W����<�o�<�-j�1FS�Ӻp��(��   (���n޺��7n���6��S�@R���      'w     �ǔJ�?����y���{[���]8Q.^P�\)j,   ����ʊn޺��wn+��B�c\����~�_2     ���      �FQ��y��sn����RI�Νׅ��466V�X    ���u��-ݼqC��zas� hYk5M��IR���      �w     pj���ɲ�G�<����]�xI�6(b, ��%I��I"�g�q��� G��Ɔn޸�[�n���2�� ��0�F����B�     3�    �i�a�7�s�u�M5�^����p��jQc�TJ�Ty�+�2e���4S��r��{?S�;9�+�3��)�3y�f��$M$/��nY�9�,��y�Ğ��<?����|f�=�"c>�y�A #�(�v�#k�@A�>��(��VQ)A�(�dm�0������	9�x_����ey�Z�A�n���4M�_R���      � w     p*DQ�������k������L�    IDAT�Μ9��/ijz��� p��i���W�&J�Di�*KS�i�4˔������駽�$���)ϳW_�E��0R���HQ=z-
C�Q�8�E��Gq�8�{-�Ǳ���^��������u��uu:�Bfc\E�wu��2     ���     N�0��y�ߓ��BQC��'t��%�;w^Q5 ��4M�������������'}%I���c���(I�{�ub-�����K��|�[|�K%��X�Ri�y��R���X��D��ky��n\����{r�2��SݿWR��      ���     N�8��q��d��_���E�Ο��KO=��ѱ"F��ɲL�nW�^O�~O�n�Qy�����{�{���zA�R)~T|/�w���rE�J��k�����AG�פ���֭��q����6�i�M����w����     8"(�    �#��w8�?˲g��99�ХKO�칳
�B�� P�z��:��zݮ:ݎ���{}�z]u�=�y6�@��8V�\Q�\�-��+�T~TU�TT�T���#kͦ�]���wn+��BfAp�Z��4M�~!     ��;     8(���<�V��p�8��u��S)b$ �.i��������;�%�NG�nW�nG�^O��AG�� T�VU)��+���j����sN�p��$�͛7t��K���*d����?I��=�6

     0 �    ��E�[��?����y�i�����ҥ�:�<��80�9��}u�]��j����vK�?O�d�1�S'�c���G'��kC�T+��+����j2��* �������_ҭ�79��� ��(�����~���      ��+�     �X���;�sߗ��B�J�ң�ڇ�9 �)�\�����;�O=����yt;���Z�j��Z��zm��^{��W�����z�Nuo�ۅ��`���Y��]I���      ��;     8���l�$?��:�\\�̉�I=��e�={NA1�)�W��w��N[;;;�z�nS`N)k�c���|�>����cE������keeY׮����E9��^����o�������^+ &     ����     ��r���Y��h��_���u�0u��y=u�i����	�SggG��m��m���w�o�~^D���R*�v����C��C{�r�����n��ׯ�ڵk�v;��g��A|,����v�����      ���     ��(���9��<��1oxdD�����.rz*�G������������vK���j�����#���#8%�0T�>���!kxx��#?� �vn�w�^z�E���23�c̏gY��2     � �    �QQ���y��s���a�Z�/,�K�5=3SD> �T�$j���i������������R�e�� �(�c��u��jdxD�z]�z]###
�`�� ��֖nܼ��׮)I�}ϳ�v� �'i��G���     �w     0Pq��9�cy���~�-�j���������R�\.""�c���kc����Mm�}lmm���: �Z�z}H###��Ȩ��wO}���i����z������y���� ��~����      O��;     �8�ߞ����y~��ySSӺ���ZX8#c���dI�<Vb�x���� ��Z��[|����F�wK�a:������^|Q�������0�Zk�/I��,      ����^     p�l�����}y�O�wX�:�._������8J�<�-�o��767����N�3�h p,��u���jdtT����;��_N�N��k�^��k/�Wl��[a�T�$?$��?!     ���%     8�Q�X���rΕ�;�^��ҥ˺x�J�}�0`�9u:mmnj���ͽ"���V!'� >;k����4<2���Q���kxdD�z}�� �s��ܹ��^�}ϳ��� ��4M�]���     |v�    ������܏�y����`��fffu��+����Q�����Z__W��������m�� p��q���q���jllL�c���v�� �N�++z�ūZ\���1.�A�m�~���"     |�    ���ʲ�ǳ,{�~g�a�/���Okhx��x I���+����+�w:�A� <!k�FGG5:6��ѱ���蘢(t4 ��N��_zQ7�_S������KA�������     <B�     &���p�}_����U��t��+�x��8."��n����[�j�����: ���u���k||\����7�˲L7o�Ћ/^���־�A�b���4M��x      �    ���Q��<Ͽ�9W����I]��Μ�1\� �ｶ���j�v��{e�"N ��z�Q�}||\cc�ށ����%]��������,k�v�?�$�J���     �V�%     O�E�������s�j+ct��Y]y�MLL��>9紹�����j����R��W �~��!���k|bb����q�Q4�X $mnn����u��M9��5�Z�Zk?�e�_��QLB     p�Pp     �K�Z�M��g�<�:�}��YQ���K�r��j��"xB�nW��u����l�j��T�烎 8����&S�
����:pj�z=]���^z�����fc\
��]�^�vA    �)@�     �&q��9��y���~_�������gt��E�aXTD �C��j�������5�`mM�Ngб  �\���Ą&&&519�j�_�[�g�y󦮾������5�� ��1�[�4�hA    �	F�     ��r���Y��D�eo��F��+�<����e	�0�����ښ����ښZ�u9� �WU.W419��Ɇ&'W��	x���ZZZ��������Ap#��������    ��;�     �eEQ��ι��|v?s�1���ӳox�&'E��
�<Sk���ֺ����\]���Πc Pc����5�h�јRc��Z�>�X���j�t���s�־Q2�;A|o�$���x     ���     >ME����<ϧ�3'B]�xQW�yVu
G�����փ�����ִ�ђ�~б  84�Zm��IM6�/�����^���הeپfYk����K�e?VP<     ppe     H��0��ιp��gN�\�姯詧.�T*��666�����ꪚ�U���A� �H	�P��55��511� 8Q�$ѵ�^ԋ/^U����,k�V�?�$�I����     �أ�    ���q�CY���9W�Ϡ�А�~��.]z��P �Z���֚j6W����$I �c����1M6�ԘlhzfFq:p"8��Ν;z�Oh{kk_���� ~5M��H�^     N)
�     �N�(�~"��ov���39�гox����e���r����j��huuUkkMeY6�X  �(�����ј����R�\t,�X�����;z��Oj}}}_���� ~%M��J����     ���3     ��pE?�e�;���~5=��57?_T6�T��\��u5�M-���Z��<� �S�^�kzfF�Ɣ���U�����Z���N�����c�ɂ ��Y��5IŤ     Gw     N�Z�6���)��?ｷO:���g���7�A��cEFN�,��l6�l������97�X  �3���jjjZS�Ӛ��V���R�����?��w��{��s�1y��eٷI����     �ȣ�    �	V�զ�����y���ۃ Ѕ�̳oP�^/2"p�i���V��j��j}����=  ��c���{E���v[��9ݼyc_��i�qA��R�􎝝��#    �#��;     '�^����<������?�"]�xI�>��*�j���{�V����e-��Wsu�� 8a�1��̌f�g5�h(�A���^���W��K/��,˞x�^��CQ���nw���     ���    �	R�Vg�$�����岮\yVO]��ɔ�k�������ZY^��ʲ�4t$  p�� Tc����YMO�httT�p�l����^}A/�xu_?;?Vtg�۽[`D     0@\Y    �(��^ѕ+���+O+�"#'J�eZ]Y���=-//k��t$  p��J%MMOkfzV333��냎IY����z��ϩ��>�c����0|W�׻]`D     0 �    8�J�ҥ<�1��/�O��V���3��ҥ�A���{�V����e-��WsuUιA�  �D�^����n�}v���|�rݼqS�=�qu:�'��Wt��0���;     �w     ���b�?�����Sl���&�=wN�p� x����/����}���*˲AG  '��V�Ɣfgg53;����AG��n�����_I�+��~E��v��F     ��;�     #�ju6I�_�����)�����gߠs��Sl���}���hy��/�W��3�H  �(��jLMifzVs��T*����^�����>�����z�9{E�?����n�n�    ��6     �@�V�������b��dCox�477Wd<�X��k}�������V�5�H  ��3�h||B�ss������Ġ#���۷���>����q��N�s���     � Pp    ���v�����ۼ��I�LMM�Mo�\MMO8v�4���}---��Ғz�ޠ#  |V�rEsss�����̬�(t$` ���s綞{����|�9���dY�I��%     E��    ��T����,{�~��FC�>�F����8V��V����tO��ߗsnБ   ^7c�&''57������:p��������cj�����X���6�K     �@��?{w^Y~���sV]m��$U�T�U���U�]���!��L`Ϙ`3!�d�$�<!d���C 0��lL�c�n���k�J�E�RR��+��;���w��{u��ޯ���������    @q���������"MM{t��1555���(҃����0���y-/-%�  �wUUUjnnѾ����$�����v�8֭[s֓'�s��eY��8n�y�$n     (,�    PR�����Olg����Ɔn�^����n�^PI'  l��o�>���Wss�|�O:	�2��~U���n�v�8ο��g$���    �\��    @�l��~9�EQ��Jcc��9�={��(j+++}J��-ݻ{Wq'�  �8˲��Р���j�ߢ]�j�N���;wt�ʥ�]t�p��A��I��W     ���;     	q]��(��(�*r�Fcc��=�={XlG��P����¼n��imm5�$  ��WUU���jinQӞ=�,��-��khhPO�<բ��mۿ`���<�    �M�,     ���y����0�����M:z츚���� ���������I:	  `�J�Rjiٯ���ڳg�l�I:	(�8�533���ZY^��:�m/9��?A��<�    ����;     [�����߆a�?�k��ݠ��#jni�gPT2���57;�۷o+����   J��ڻw�Z���Ҳ_��%��]Ǻ57���+O���8�#�q~:��|,�y     �M��    @������oczs�FMM��9�ֶ�|�EcccC�o/��  � �q�w�^57�W���J�RI'yE�fgg4|uH+++9_�q�[��}}�/�     ��     ��yg�8��1�P�ר��ё�����b;J���n��j�֜>x�8��N  ��,�RӞ=j�ߦ���U^^�t�7Qj||\ׯ�(�N�|�u�ڶ���Lf8�y     ��Xp     �*++�lll��1�\�Q]�KG�U[[�,��w����%ݚ�խ[sz��Q�9   x�eiwC�Z[���ڦ�������C���Q]�6�L&��5,˒�8�<���t:=��D     v4��    �?U����1�G�8�s�@EE���������v����E���ja�K�   �XMM�Z����ѩ����s��f���訮]V9]ò��q��c�����    �3�    ���z��KƘ�����������?����vN��@Qy����n���ܬVVV��  @�544�����Q���u�ڈ��FEQNװ,˸���A��$��B     v�    x
���\E�sE�����ý}:t���w��ܿ���ݺ5�����s   �EXvG�X[[�իW5=5�8�s��m۫�m��1���s     ;�     ����EQ��a��2�8��{z��Deee������f�f5=5�I�   P}}�::���֦T*���[ZZҵk#����y��q�G���L&��y�    ���    @R�Ի� ��0l�e޶muvu�ȑc*/g����,��LOkyy)�   !˲��Рֶv��w��^lKO�<���U����|�q&|���t:}.�i     �4�    ؄T*�e���1�l.�e���]G�WUUU��[^Z���ffg����t   ��q�o_���;���"�q�N�r��]^����|�u=����tz.�i     �$�    xk����1�G�8�s�@ss��?��ں|�����ٙi��L����I�   �����-���ޡ�{�ʶs��17;���+Z^^�i޲��q��c~X�J~�     (,�    �&|��Ec�E������8qR��M�N
&����ܜ���t��=�q�t   JTYY������ѩ����s�M��H��������a�v�q�A�/�    @I`�    �o�y�?��W�(��e��z��;�ֶ�|�E��ܾ�ٹY���*M�I   �a***��Ѯ��nUW�J:x[�����ڵaA��5l�^t���w�[    ��Ƃ;     _�y��(�>�aW.�eee:|�O��m;���*�c=|�@�s�������F�I   �$���^�]jkkW*�J:xK�q�n޸�(�r���8�|���t:��<�    �-��    ��R�T�1��1gs�w]W�����O���;ȫ��EMMOjfzZkkkI�    oʶm��׬��N57��q�#1���Ғ�����\��p]���y�y:���c     ��    ����u�����q��=�eY���ё�G�J��ȋ����LkzjJ�=L:   Ț��jmmSgg����ԃ4x��߿�ӼeY����'$��    `{`�    �#���/�(��(�rz����{u��jkk��EǺw���'�4떢(J:	   ȋ��J�w�����*��������y]�|Q+��9�۶���/d2��-�i     =�    ;JYY�wc�}��s���Р�'O���Q�=|���)��Lkcc#�   �`,�Ҟ={��٥���r'�$��DQ���Q�_U&�������<�������<     ��    �!�J�c��s6����J?~Rm���N�Z:���Ԥ�������t   ��<�S[[�:;�����Q\2��F��jll4�k��;�y������<�    PtXp    �:��c>Ǳ���y��;���q �JEZX����n/,(�㤓   ��P]]���.utv���"��V��58xEss�9�[����� �')�#�    �Xp    �,�u��(���(�R��Z����N�8qR�T��@�,--ijjBS��Z__O:   (Z�e�i��tP��������Çt��%=�?�y۶���� >��4     ��    ���J����a�7��={��������;�I������Iݽs'�   `��}_�mm:p��z(s���������Ǚ�}����syN     Q,�    JFuuuC:���1�\�kjju��)�ݻ/�i@N�ݻ���	���*M�9   @IhllRww�Z���8n�9���0����6"9]�uݗ�1��8�u ��     IDAT    $�w    @I�}�� �Wqg���J�t��quuw˲�UF����5=5���	-//%�   �,����ѡ�����'��.�Nkh芦���q��e����v?U�<     �O�    �ZYY���EQ�;�Y۶u��a����y��6%�cݽ{G��ukNQ%�   �(uuu��9�����"A�>ԥK�������y�8Ώg2�O�9    �-Â;    `[J�R�ƘOc��2�g�^�:�]55�N6m}=���)ML�iee%�   `�s=O�����9��:NuGr��u��y����4���yߛN���    @���    �nl��~��8��l��w��ɓjnn.D��8ֽ�w5>1��[�8�   (R�����>������tv�04�9����2�d=oYV��A�㒲�      	a�    �mx���0�]EU������G����AY���z�tZ������>    [��<utv���G55�I�`Z[[Օ+�5;3�Ӽm۫���l���4     
�'�    ������0?�aw���e���A=zL��"xK������(��   %���Q==���&�q���s��}]�tA�=�i�u�k��|����x��     �+�    ���<��Ƙ�q��=�޽�t�Ԁv���xS�LF��S���R�9    򬬬L]����9���ʤs���q���I^���F��eŎ�|��ÒL�    xz,�    ����?j���(���������Sji�_�4�M=z�H�㣚��Q�'    �:˲��ܬ���o߾�s��d2_��ب�8�z޶�5�q>���    ��Â;    ���R�Nc̟c�g;�8����t���W�c˄a�ٙ�����ÇI�    HHuu�zTgg�|�O:;ē'Ot��yݿw/�y�u�\�������<�    �3�    ���<�׍1����v���E�N�VeU��9I�Ӛ����͜^   �49��ֶv>|X��uI�`�X��ׅ絶����eY�뺿�?��    ���    H���?d���(�����޵K��w/���ָ{�F�nja~>���   �9�t��A���*�����@V�1���7o(���S�m{�u��g2�O     �Mc�    �����}�L�SƘ�lg�Uo_����d�N!�o0�hfzZcc7��ɓ�s    l3�T�zЁUVV�tJ���._�������]��}�{���n�9    �Ma�    ���~����8������>����B�߰�����qM��+��$�   `��m[m�:|��jk��A�[����K������eY��y���d�U�     xK,�    �T*��� >�aC�����:5pFMMM�H�aaaAc�7u�vn��   ��iڳGRK�~Y�mQa�ڵ]�6�(���w���?�N��V�<     �-~)    l�
�u?���q�ՠ�:�ۧ��~�v���E�fggu�ڈ��   �CTVU�����{z��~�9(Q+++�x�|��v]�ec��JZ�o     �    ���<���W�(*�v���]'O�RyyE!� ���illT�c�d2I�    ء\�Ugg�:���]I�D�����J��Y�ڶ��8�?��
�    �7��    (�T*�i��3c��lg���50pZ��5"��Ǐt��M��L���v    (˲Դg�<�斖�sP��1�q㺮��t?���ߵ��>S�<     Xp    ��y�b���8��l��Qo_�z{��8N��C�q���9zCw��I:    �R]]��U[[�l;��k�m=y�D.����g=kYV��oA�SH    �p,�    �*�J�+���qE���mnn֩�3���*Dv� 491��ћZ]]M:    �RQQ������G��%��391��������zֶ퇾��������    ءXp    �K��n�yg�����:~�:::хl}=���q�޼�L&�t    <����խC����2���L&�����8���w]��Ƙ i=�u    ���w    �S�<�a��(�ʲ��m[֑#G�n��=y�X7�_��쌢(J:    �ʲ,����po���~��<����Г'O���m{�q����w�    �AXp    䬺��!�N�s6�ٺ�z�y�Y���";ԃ��u������N   �-��ب��~5��$��Ǳ��F54xEƘ��]�,++����ջ�    � ,�    r����A��8���u��t��q8pP��m)�^E��uKׯ_ӣG��   �D����po���;��F^�����}{!�Y˲��y�:�����    J�l     ���~_��
ð+����6�8����B�a�	�@�c�y��鵤s    �(TVV���^uuw�q��O:�m��L��Z__�z�q�[��{ccc� i    �ł;    `�<��c���qlg3W^^�S����V�4� ����d2I�    @Q*++Ӂ��t��A���%��m.��hx���Fo*��f-ˊ\��� ~�@y    �Â;    �m�R���d2E��l�,�RWw�N�8%��
��buuU7o�������$�    ۂm�jk�P�UWW'��m����:�u-..f=�8�=���?�N�+@    ����    x+��b��{������3Ϫ���]�A�<y���F4;;��)q    ��fY��;:��ק]�j���6E��_ѵk#
�0�Y˲b�u�8�,)�a    ����;    ���}���1�EQU6s�����:x�,��N������~mD�I�    @ɰ,K�������?��,//����u��ݬgm�^�<�766>[�4    �6Ǧ    �[�\��Sc��d;�o_�N�yF�������0?�k�G�����S    ����׬��~566%��mlrbBW�\R&��z�u��c~@R��    ��ł;    �|��Ac��EQ�Ն���:~���{z
��Ǳn/,hx��=z�t    �(������WsKK�)ئ��Ӻx���f���m{��������    �!�    �T���s9����Mg�J�
хǱn�����!---&�    ;Zmm������C�ţddoa~^.������g]�}��ݒV�_    �N�U    v8����;QUd3WQQ��g�Qs3��!{QijrRׯ�hee%�    �߲��F}}�,�#'�LFW._���Dֳ�m�����L�
�    �&�5    v�Z�u?a�y)����8qJ���%,�BMMNid�jN��    �NeU��z����͢;�v��=����Z^^�z�u�sƘ�D�r��     Ŏ_!    `�<�a�ZEe��UUW�3ϪiϞB��Dc499���F�N���    d���R�����G��$��m$C�����8�Y۶���� ~�@y    �"ł;    �,���~�s6�!۶��ׯ��~d#+Aht��n޸�L&�t    �)TVU���_��]�m;�l#�>�o�ӓ'O���4w    �yXp   ����l���(�R������ٳϩ���Pi(A,�   @骬�To_����YtǦEQ�k�FtmdXQe5k����?��d��@y    �";    ��
�u?n���l�l�֡Çu��qVcӌ1���#,�   @�������>uw��qx�6gq�^?wN�=�z�맹�G�j��     łw    (a����1�#QUd3W_�[Ϟ=����B���A�ћ7t���   `����P_�uus�;6'�"]�~M#�Ws=���f2�?.P     a,�   @iJ�����ڎB��v    �ߨ�����^���ȶ9�ooqqQ��{-��ܿh��^I�     %�w    (1���1�QUf3�{w��}��v��*%��nrb;    �ۨ��ґ#G���)��4�ZǺ~mDù���y�oll|�@y    ��k    ��uݏc�~6C���ȑc:���Cg��04���е�a���'�    (b�UU���WWw7�9�m--.���_�Ç9���c��I2�/    l5~E    �PVV��A|<���l��̳�i׮]�JC���HS��R:�N:    ��쪩Q__���;Xt�[��Xcc��rEa�ݮ�m�O����^:�~�@y    �-¯    ��Y����1��qo��q=v\���2�RE�������֒�    lcuuu:r��ZZ�'��"�����ϝ�Ç���,+v]��A��@i    �-�    lS��	���a��f���Ng�{N��u�JC	��X���48tE+��I�     J��ݻu��	�ٳ7��8�u��u]�:�(���u��8��d2#�    �    �y���Ƙ�ͩ�e�po��=.۶��m�oۇ�����t    ��566���jllJ:ElqqQ�^��?~�՜eY��y�{&���J    �    ������A�cLo6s555:��󪫫/TJ��;wt��%=~�8�    ��g�^�<y����M=�iT����ջ�    ��    �Mx��ύ1�Ǳ�ٙ�xj�1ٶS�<lc����ݻw/�    �eY������񓪪�J:E��Çz��״���[�,�2���7A�Z��     yĂ;    �Z�u?c�9��PUU��=���ƛZ\|��᫚��M:     I�m����ґ#�T^^�t�P�ҍ���qV���3�|�����    �w    (b�����(�6�Dײ,<xHǎ���pj;����e]���L�)     |[�����C:��'����A�w�^?��VWW���m{�u���d>V�4    �Sb�    ����Ǎ1��f���RϞ}^MM�ڎ�+�^���UMNLd}�     I�}_��Gt��A�6��73A�˗/ibb<�Y�u?�������    ��    Pd|�?��_�aؐ�\Gg�N��B�a��d2�vmDc�7�<�    l?���:z���;dY<��7[XX���������l�~�8�{� �R�4    @��   �"����	��_�q���5��50pF�,�vE��&'54tEI�     ��v����cjmkK:Ef}}]��{M�o/d5gYV�y����d���    �Ă;    �z�u�d�9����}���ϩ���P]؆�8�����������t     y�g�^�8qRuu�I����q��+�u����g]�+//~yy�A�     Y`�    �y�?	���������8:q�<T�4lC�o�����z��q�)     \{{��;�ʪ��SPD���t��y�q�՜m���?���a��     ���;    $�q]�cƘ�f3T__���=�]�j
Յm���G�r���޽�t
     [ʶm�8���#*++K:EbzzJ��{-�%wIr]�3Ƙ�d�_    x;,�   @<�;��g�(����eY���ב#Ge�v!󰍬��hhhP��39=�    �T�����~<tH��$��"�4K��<�m��� �T�4    �[�    ���y�j���8�S������w������e�_eH�LFCC�:w�kz��q�9     $.CݹsG�3�*//WMMm�IHXmm�\�ѝ;ٿ�.���8�?������    xlE    �֩w]�KƘ��uvvi`�\�+T��(�4>6����d2I�     P�v74���544$�����uML��<�8�d��Hz��*    ��a�    �@YY��A�GQm��v��t��3j��(`���w��ҥZ\\L:    �m���E'O�VUUU�)HH����?�Ǐ�|۶7\���L&�gyL    |,�   @�y��A�d63��M:��󪬬,T��Ǐ��K�w�n�)     lK�m���C��?"����A������~ZƘ����f���<e    ��   �@���[3�̫a�nvƲ,�9���#�,n�v�t:���!MNL(��s     ��|�Woo�>$�v����yC�.]|��8�3�yދ����O_    �VlK    @x��Ƙ�;�cw�3UUUz������i��1�~��n\��0|�S�     ��U�k�N�<��斤S���8�>�9=z��eY�q]�CA�f�     �    �_��n��O�������3�<�P]��8��Ԕ���(�N'�    @�۷�Y'O�Ү]5I�`�<|�@_����v=�u_6ƼG�    @���    y�yމ0�EQ]38}F��L�6���C]�tA<H:    �Ų,uuw�ر*++K:[��W^���[y���8�l�~wW�vQ    ����    �����Ƙ��q\�ٙ��F���VSSS!�P����t���t���֒�    `Gz�葦&'乞���eY�W�jjj5>>����q\��O���Eѫy�0    �Pܕ   ��I���Yc�K�<tX'N��mۅ�B��P�7oj�ڰL$�     �n׮]:yj@��5'����/Iw����u]׽h�yQ�z�/    ;�    �#����QUov���\g�{^{��-d���쌮\����դS     ��ؿ�U'N�RUUU�)(���y}��*ȵm�^t�A\.�    @�s�    �����_4��n�e��ٷ�Y/}�T[[[�4�Ǐ�k�~U7o\W���     ���%���ɄF�����TUUkrb\Ƙ�_;��T��}?��    �8Np   ��\���1��ض�cǎ�po_!�P����uuhP����8�     ����
�8yR��I� �._���7o�;\׽h�yQ�zA�    J�    �I�����QUov���J�?��v�n(d�T����!e2��s     �Sjjjҩ�3���D<�__����=�m/:��� .��    �8I    �v���/c~7�����om�K/�S�՛އG	��^y�eMMM*äs     @���jbb\+++jll��I'�)�WTh��EQT���8��}ߏ�0�JA�    J '�   �[K���Ec��pG�N�VwOO!�P��鴮\�����S     @���������e��}�z�+/k~�֖}�뺃Ƙ�$���K   `��.    �Dyy�����r�3�v��_TM���i�(����	��s     �ٽ{�Ψ~��S����F48xeK�Ӷ�'��|g�[��    �M8I    @1r]���#q�mv���S����TQQQ�4�;wn땯��������     �t:���	������Q��&��,jfzjK�3��T�?�n:���m�   �6�	�    ��l�u���=�pGg���]�.���U]�|Q���N     E��};~B��=�,�o�tZ��ğ&����l�y�$�X    �   �����A�(�6�>���]z��U[[W�4�(�4>>���+2�g�     ��������3ڽ�!�l�����ab��8�]��[__�ڣ�   �H9I    @1�<�}A|>�����om�K/�S����LC���^��_izjJQ%�     ���zZS��ZYYQcc�\�M:	oajrB�L&���*�y�7Eѕ�B    �Hp�;   ���A�c����8:yj@==
��"����+�/iz���     ��R�:y��;:�N����>�$�!I�< �GIw    @�Xp   �cUVV�Y__#ö,f�����ݻ��"Ǳff�u��Emll$�     ��Ʀ&�>��jjj�N�����Rw��I:�Ǚ���xvyy�8��   `�9I    @��ʾgcc�\E��Tomk�K��.UUU2E��Ç��+_��ب�0L:     lck����W�jhl�m�I'����f����t�7�q\4�f    IDATg���|�?��D�=    ��Xp   ��x��kA�_q����m�:uj@'N���p�d2]�|Q.�W:��t     (q�������VUU�v�ڕt$MOMie�x�%)�c7���}�,ÿL�    ���t     l���_6Ɯ��@EE�^x����P�.���i]�tQ���I�     ����U�U^^�tʎ������ݻ�tƛr]��1�%I��[    `+l�B    ��|�?��׌1u��ٳw���E���2EbeeE.��;�o'�     v�[ss�{玎;��eY�Q�� 0I'�%c�Y�q�:��B&���t    ��t     ��y�3�|.����������g�����RǱ��F��W_���R�9     `���H�o/ha�����9�=�W�dLq/��q����=ϛ���J�=    PH,�   (i��}$���do��z��u��!N��?~�W��&''EQ�9     `[__���2���dۛ�9O)�Bn�}q;���<�#��O&    �¶   �RU���ƘC�����/~����
م"���h||Lq'�     �M*��t����לtJ�[Z\ԧ?�Igd�u��Ƙg$�$�    �Ƃ;   ���y�3a~)�����ttv�̙3r��i(��p����%�     �ZZZ4p�UTT$�R����t%��۶W�yg�n   �|r�    �|�<�g�1��l3�wGg�<��ǎ��������^{U��WA�9      okyyYSS����T__�tNI���҃���I�~�p]w%��ג�   �|�w    ��v]��Ƙ���@ee�^|�w������,�c���jphP��v     �M55��3�<����SJ��?�=z�(錧��Ǎ1?�t    ��    J�n�q.�aؾف��&=��;�J�
م��,/����ݻI�      <5�q��ׯ��~�F��ğ���8N:%/Ǚ�p@����   ����   `[�<�0�EQ�fgz��t��	Y�D�*�"]�6���aEQ�t     @^�����3gUWW�tʶ633�׾�j�ye��ZYYٻ�����[     WN�    �+��>d���8���|�u]=��:x�0��%����z�+/kff�dN�     ����&'ƕ�d����i�9�����3�*�c/�����Q]H�    r�F   �m��A�c��|uu�^|�K���)dd���Р�Fo��     v��]���3Ϫ��)�meccC��ğ����<��� ޟt    d�w    ��.�u�cnv���Yg�{A����ޱݻwO��8Wr'n     lVGg�N��7�M�vmDC�W��(8�u�cNKZK�    6�w    ۆ��G�1_��h�f>oY���U�Y�?�(���ҥ����L:      q:}�57�$�RԢ(�_|�Z[�;߶m/���|&�I�    6�I:     6���	��q�o����ޡ���K���-}��/����I�      � 433���U55����LOOizj*�-�qYE?�y�TECI�    ���n   @��<��A����|���F�|�{���P�2$accC��x]CC�2�$�     Pt�<y���)UW�Ү]�z�E�^��+
� 锭fGQ�^���EQ�I�    �[�C    ��w]��1��fZZ��瞗�y��BBn���7����t
     ����ѩS���~�)E����|�b��r]�Uc�K�¤[    ��a�   @Q���ط��q9�=�����ӱc'dY�ꔚL&���˚O:     `�I�R8}F��mI�$*�N���ߧv�����8�|�?�N��n   �o��   ���J�ޕ�d>EQ�f>ﺮ�}�9����t�jvvF/����F�)      �Z{{�N�VY٦~v+9_}�+�uk.錢a��zYY�{����I�    ���$     ��y
��?�q�m�󕕕z�ޭ={�:[l}}]��{M#�W��-     �i-.>��Ԥ*��TSS�tΖ��׍�ג�(*q�a���y��(z=�    ���   �hx��� ~l��ojj�/~ǎ=q������78�     �@���5p�̎�mmqqQ���g�&锢�y�oA���;    @b�   @q(s]�Uc��f�{z40pF�m�[,��hp�&�ǓN     (y�TJ��<���[�N)���}�����r�)E�u�Ac�IA�-    v6�   $*�JuAp>���|޶m�QwOO�Ӱ��u��וN��N   ����;�������yΪ꫺���g�\.�$w�%�K���+�Nr	�ȀcAN ���%F��P� 9Hq�(Nl�I)��H�Krf83�px/�<�������9�G�49�]3]UOu���������b����- 8V��^=����8N�Q�*C���i}}-�(G�eY��>^�V��   ����    1�T�|��gQ��׳ϞQ~l����F����7_gj;     @�2�����S���J:JSDQ��/_���B�Q��4�����Z�GIg   p<YI    p<���{���q�v#�sz��?�`.��hh���e���ZYYI:
     ���n��T�z]ccc2M3�Hw-C]�tQ���IG9��8��0����lEQ�J�y    ?Lp   �v���#���j��'&&�̳�u�W$ga��w��O�_q'      ���ק�O=��|>�(w�^���Z[[M:JWp��}��'�   ��B�   @;��m_	���F�=�G����/�b}}M�\��R��t      |�0���w��L�h|9��֖._zI;;;IG�*�m���$Ig   p<�   ����c�Z��0�Yo���|�)����VGC�DQ�w�}G����     ���z��3��rIG�Z���x���0L:JW�,k!�G%��   ��Qp   �r��<��(�zY�N��ܙ�mu4���vQW�\���F�Q      p�L�Է|H?�mYVgMs/�˺��u-..$�뙦Y�,�Y���L:   ��F�   @K�������q7�����Μ=����VGC�|��z��7��     p���������t�Q��>�����wA�q��0B�q���y�$�,    �w    -���y��nt��Դ�~�Yٶ��Xh�j��W�]���R�Q      �D##���#�hll��gGQ�O>�D?y�]U�����0��q���y��I:   ��D�   @Kض�gA�j��|�!=��we�L�s���~�y��t      �H.����K'N��e�vhE�Z��>�H��j�ZK�Bcl���� ����   ���   �li۶_���F�����)�sｭ΅6�}_7^��O?�y�Q      �&�mkzzF3'Nh,?&�q��o�R��Ңn��Tk����)��yl�~?��%q�   ����   �i���)��_�0��z�u�ܙ����Zm����W�]Q�\N:
      b�FFF422��\N��9���ɲ���{�z];;;������VWW���ݦ�8˲V���#�ry%�,    �w    M�8��0_��(�����>�;wA������H��~��{L�     �/�J��J�eۖ,�VG��H��Z�)��#�LӬY�u���W��   ���   ��\��W}��'q��=�##:s��醺��`�]�zE��kIG      � �0B�q�u������    8�*�    �Wq]�w}���8��F�Ϝ8�3g��u�VGC�}���u�����t       �3�(�5۶kQ��t    G�   �5�q�����������{�q/E�2�����Wu��IG      Ё��c���F�9    M�J    �Ӷ�Ap��Ŧ�'�|J�չ�b���z�e���      �kض�rg$�Ig   p�Pp   p�,�z;Ó�,v]W�=wV���V�B�q����]���w�|      �`�e}�ᣒ*Ig   ptPp   аt:}��y�GQ�md}__�Ξ�����VGC��e]�����֒�      ���,k�u��V�չ��    8(�   hH:�>�y��E�������9{^�T����B�~�s���u��t       G�i�5˲.��-�,    :w    r�7� ��8��F�OO���g��e٭��	�Po���>��IG      ����5������    �lV�    t6۶'�?h��~���ɧN�4y�qT�E����0�t       �Ì��ض]���J�a    t.&�   �J�����������#������Hh�O?�������0H:
      �.�8�����I�    Й(�   ��l��� ~����i���gt���V�B����믾��ٛIG      pض�σ �KI�    �y(�   �"۶��A|��Ů��̙s��[�-R(t��e���$  �-lۖd��������ÐeY_�ò,�����q�0���0����
���A )޻   ��m�oA�=I<�   ���;   ���,��0gY��קs�.h``�չ�"~���|�uEQ�t  �}�iʶmY�-۶eۖlۑm[�,[��[N����¹eY2MS�y�������"�c�a�(�E��ax�q�W�����A�v��� T�{�����   Q�e͆a�mI���    �G�|    M�N�Oy��fE�F����J�ӭ����j�v�������  ���8rw���r�na��B���"�e�2ͯ�����-����[�[�����}���w�'   ]���M�u�V��Ig   �<
�    �8�ca^�������Ԕ�~�9ٶ��hh���U]�rY�j5�(  �ٝ��(�r庩�Rz*��뺲mG��*�J�q�#;)w.y^]��?���������8N:2   :�i�5˲��}�F�Y    $�O   �c.�J���yǱ���{�WO>y�������7^WEIG  �0��R�릔J}vsW���v����8ޟ �y�<ϓ��U���<��Z�N  ��2#p]�W�����t    ��	   �s��
�࿉㸡�>��}��V�B��u]�zEKK�IG  m�����t�sE��	�LZ�T��::V�V��%x��T��U����V�)äc  ��Èl��������    H�\    ǔ����y�Q#k��O|_�}󛭎�(
���%��夣  �&�mG�LZ�tF�tZ�L�)��$h9��T�{{�k��j�ժ��j�V�
� �   ��aĎ����y?�,    ڏ�;   p9��G���V#kM��駟щ'[-����7^WEIG  w�0�R��{&�[d��ض�#/�"y^]��n�Z����劢�	�   ��q�����7�    ڋ�;   p�ض��A��Fֺ��3g�i4�ou,4Y�^�+׮hqq1�(  �k8���)��R)o�6[��Xa(�b���a(�o�٭��EQ�$m��L�����^�p��C��/_�`Y�{X�-�0����8V�^�m����{�Z���IG  �$�q����_O:   ����   ��0m��q�Y�������f[�M����+/_V�RI:
  ��$�t:���e2=���QOO�zzz(-� ��0�{�?�p���YY=TG
�PQ)�n=���걂 �xvg3dۖ��\ޒi�2�ݟ��o�J��-�ڻ�e۷n����eA�R)�R�|�VV�VS��+    �R�m_���s    h
�   ���ڶ�V�jd��@V�/\POOo�s��~��Ǻq㺢(J:
  ǎm۟+�Vd�d2�n{��}�����ϕՃ/��/�ٿ<%�w���Y��B����8rw��9����T�V�P|߽��)�   h۶�	��qI<�   ���z�   8�,�z/éF��J�R�΅&
�@��zM�7o& ���J��Pb�-����t���y�J����?{���p|�*�;�+׽�����~�{��&���*�����&�W*�����  t˲��0|XR)�,    Z�{�E   �L&3U��߉�(�����)=��s�,����D��ۺ|颶��IG ��X����^������oﾷ��+�NZ�T���yu�뻷[�w��
�q�q�����TJ��R*�R*�V*����U7}������e���hggG�JYa&  �ȱ,k3�J=\�T���   �5���a    �q]��A�EQ����Nݣ'�:-�4[M�0?�k׮0% �Crݔ�����ӣ�����G�-�8�������j��<��+�{򼺪՚�����::�m��d2r������{:��+§eYV�1��<�J%��T.�U��U.W�%   _�4Ͳ�8O�����   ����3    �R:�>�yޏ�(rY���ǟ�a�ᨈ�Xo����､�  p��Ne�Soo���j���՚j��j���[Sع ǁ��S�����2����X�ߝ�^V��;����w��  ��4ͺeYO���F�Y    4�   �ˤR���y�?�㸡&ǃ=�G}�ձ�D�ZMW�����夣  ���Q������}�d�:*o��q�7}��Wd�~�qM��%�x�&�V|O+��(�ٝT�=�bU�5���hggw���vIA��,  �x3#H�R�V��(�,    �稼s   ����k����8�̓���'��}�w�7�M����+W.�Z�& ��bY�~���}:�N:ց�0T�z��^�B���8���t-�0����/M����4;�{�ZU�TR���Ri��Τw  p��9�����i�Y    4w   �K8��A��q�<�4M�~��8q���$?���z��7�q�Q  H�a���Q__��٬�٬zzz��owA�r��J��j��J��r��Z�&���@'�m[������ݿ�U��d�ZU�bq��^*�E\,  ��a�m�����>�,    �s?�   �0۶'��op��}�&&&[M�^}�fgo& ���|������4����X�zM�jM�Jy��^��NY��%@�ض�?�}��޳��S�m�V+{��)� ��eFlY����?O:   �á�   q���=��~���:{�FFF[M�S*������J:
  mẩ����������h����+���Պ��j�*ߴc�a(�ɨ�g���٭W�e%�6QjggG���*���.��  t�u�S���äs    �{�  �#�q�?�}��Y��dt��488��Xh���E]��2E @WK�3���l6���ޤ#���<�J����;;%��I�4�uS���WOO�z{{�w��4��X��/��J;��:  pT9�����I�    pw:�S    w�q�����_odm��_x^���U�W�ɻ���w�a
, �������>���+��jp0'�q��%iw*{�RQ�R�/����������R�e�Ox���W__����:f�{������vq��EQұ   �8�����o$�   ����   A�m��A��F�d��p�ye2�V�B��k�\���\�Q  84�u��?�l6�������e�fұ����u��8�����Wx/jkkK�ϷM ��f��?��_J:   �;C�   8ZL۶_���F���J�R�΅&(mo����.�� �]���Q6;�_hO��X�JU�ҶJ��J�����a�p. �3�e���W}}�P_߭�{��Պ���	�[�V�IG  �۶/Ap.�    G�   8:L۶_���F��c:{��l�iu.4��ܬ^y��O:
  s]W��r������J��sk2���n�}{�(�߭ ��eY���S__�����&��&���<�[������j�Z�y   n�m����1|u   pPp   ���?�    IDAT��w� �f#�'&&�ܙ��,�չ�����~�M�1��  :����l6�"�����}/�< �	l�Voo���f���/�u�S�UU,U,��QP�^O,  �m����	��   ��Qp   :�kY��a�����i=��s2M��.]�zE��sIG ��,K��48�S"9�0��Ny�̾�SR�\N$ 5��ڟ���ׯ��9	}�W�Vݛ��M�e  ��eY�a��$��   :w   ���Y��A���,>y�N�~F��S�N����K_T�XL:
  �,���`V��9���׫$�B�T������V�m�  ݬ��go�{VY���$�"��Ύ���������-�a�@  p�X�5��$�b   �P�^   ��5�Wn�7������'��}��G���._��z��t �1g��٬r�����v?���H�RI�▶��*�L��vr��{�L�lk�8�U*mkkkK��*��㸭  ��aY�J�Hb	   Ёh�    ���o�R��4���F�?��Cz���ZM�?֍�EQ�Q  ǔ���4<<�\nH�m���0��]�+�o�X,�{ :�a����/���8N[3�a���m
�*�U���z>  �~�e���7��   �v�  ����3Y��ދ�(��z��GC�z��u}��ϒ� 8f�������G����S�VU�XT��[j/�Jm= ��tF�lv�������k��677U(�����Q  �)L���d2���夳    �w   �����S��EQ_#��{���Z�T�Vu��E�ד� 8&2��r�!+��iZm:9��NY[[����}�o�� �vr]��	�}}��m�0������ml��  �4��T*�P�Z]H:   �]�  ���A܈�(s�Z�0��������f;��
��._zI�j5�( �.f���٬r���Oi�5QwssS[[����r��{R��66

ðmg ��`���ߩ�j�&�    w   �#����^�=}�Z�0��O�{�юh8���Y]�vUa$ Ѕzzz�&�ippP�i���j����MmmmikkS���\ ���)�r��ip0�t����ME�m�ݹ�  4�4ͪ�8߭��&�   8�(�   	s]��r{꠵�a��O�ԩ{����{�魷�H: ���������FGG���ۖS=�S���7wC�Z�-� �����m$���!�R�)��jU

����R�m9  M��  ��@�   H���	��z#�v�4��3�jf�D;��.�a�W_���7?M:
 ����l6�Wj��uݖ������6U,��]T�Tj�� ��'��(����]���Ň���66
*
��((Ö�	  ��4k�m?�y�{Ig   �+
�   @B���̳�izz��p��ժ.]|I���  �0�q444����4���E���-mllhssC�r��� �e���z��ihhH�lV�a���0����Ba]�BAA��<  p����Y�����o%�   8�(�   	p��0�FQt�V˲u��Y��O�#����.]|Q�J%�( �#(�NkxxD��#�a��m�Z����mnnjccCa��<  �iZ�f�7��閞Ǳ������뼮  ��K�O���f�Y   �ㆂ;   �f����bE�Akm�֙��466ގh�Ks���v�*�@ ������h^CC����o�Y�Sڋ�����֦J�RK� ����r����G���d����^��U(T(��X,��,  ���J�O���z�Y   �㄂;   �F����b���Ϟ;�|~��p���=������8�( �g�sٝF�J�Zz^�Z��Ɔ66
���RE-= �v0MK�ܠ�����)�ɴ��z�������[[[�� ���   �w   �M2��ӵZ�F������hxx��p�0еkW57;�t @G3��ht4��Ѽ\�m�I���^(��R���,  :ŭ��\NCCò,�eg��B����5ml(� p���۶}���kIg   �
�   @��/�ql��q���<��V��u��KZ_[K:
 ���lvP�����q���U�U
����P�Ȕv ��f��w���(�N��,�󴾾���U�EI�� �v�a��e���j�Y   �nG�   h�t:}�^��y#�v&�w�b���/��r��t @Giߤ�J����5
�*�J-; �����w���f[v�����(heeY��[�� @�ڛ������&�   �f�  �r�t�(�w���e���%y��t @G�|�}T��j�)qk{{[kk�Z__S�^o�9  t3�q544��Ѽ��r2�%���u���im��dw  �m�J�g}߿�t   �[Qp   Zd��~1�c砵�����h�r{��䓟��*����  ��۫�Ѽ��ƔNgZrF������ڪ
�uAВs  8�,���`N����mxM�]�� @�2Mӷ,����'�   �F�  �p�� .Sn�����}��c  40pkR{^�Tk&���5����PX��֖�8n�9  �3�ajppP###i���Z����U����T*��  �^�iz�e=����Ig   �w   ���y,�W�(��~ąa�W^��ٛ7�� H@*�V>���Ĥ2��Lj�T�*
*֙�
 @��M-CC����o����KK��V�-9  ��^��I���J:   �M(�   M�8�w����Ak]���?����NT��u��KZ[[K:
 ��l�Q>���ؘ�-9c{{[kk�Z__S�Vk�  ����FGG5::������Q,nieeEkk�
��%g  �֢�   4w   �I\�}8�Q�}�TJ�/<�\.׎h�C�bQ_zA�r9�( �60MS���^�-/�4�~F�R��ښVV���
 ��J�522��Ѽ���_E�677������u�q��3  @똦Y�m�q���K:   �(�   Mp'�v&�w�Օ]�|Q��% �b���W>?&�q���g��U����  ��N�5<ܺ�{Z[[��ʲ��b��  �a�f�q�G����Ig   �:
�   �!���`oPn?���fu���a�t @��Ri��yMLL*��4}�[����U*�� �v�.��j5���jii�o� �0M��Wr�(�,   �QF�   8�;)�;�����0��N����o(�㤣  �̶m�hll\�\���Sj  �ge���q���7}�R����e��������  ��4͊��j�O��   U�  ����dN�����(�9h��8:�iG4܁8�������G|k, t�04<<���	�0̦�_��������UJ�  �Kz{{5:���h^==�mpG�(R�P��ʲ66
\� @2M��J��V�sIg   �"
�   �]�d2��z��Q��ֲl�?A��|;��A��W.kaa!�( �&�d2�����\�m�޵ZM++�Z[[U�\n��  �{���)��kllL�T��{��u��,kiiQ�Z��{ ��1M���d�Y.�W��   5�  �;���?R.�?��({�Z˲u��y����w�V���K/ic��t �!�����MLL*��5u� T(�keeY���M�  7������Ϗ�q�&��X���ʲVV�EQ�  w˲��0�ě
   ���   ܙ�i��DQ4t�B˲t��y����#��N���^zA�R)�( �C���ٟ��̂X������ʲ����a��  �v/���466���QF�>��@kk�Z\\���N��  w�4�BE�J�N:   pTPp   �gY���0���4M=w�&'�ڑw�����_T�^O:
 �.�rZ{�R�����S��7  �W�mG���W6{���ݑR����E���p�  	�,kqo�{5�,   �Q@�   hLz��>y�B�4��sg55E���,���ʕ�|� GP�&&&�Ϗɲ���[�׵�����%U*���  p7zzz�ϏillL�t�i��a���5��,kss�i� ��Y�5�Wrg�
   p 
�   ��\˲>���AM�ԳϞ���t;r�������W_Q�IG 4ȶm���599�������
�u
^  ���f4:�W>?&�q���o�Y^^���M�  ̲���0|PR�t   ��Qp   ��i��{A<p�B�0�̳�if�D;r������ɻ�$ Р���&&&422*�4��g���(heeY�BAQ5e_  �V3MS###���544$�h��{QimmMKK�*���'  8��gߖ�4   �+Pp   ��i���A<|�B�0t��3:y�Tb�Qq��k����% p ˲466���)���6m�J����E��,3�  y��jll\�dz��o�\���VV��a��  ��m�oA�X�9   �NE�   �
�m����������o�:�@��z���f�� ��LF�����m�M�3�"
�ZZZ���fS�  �4������T>?&˲��gZ]]��¼��rS�  ��mۗ� 8�t   �Qp   ~۶_j���~�1}���Z	w��<]�����V�� ���r�������p�v�T�Z^^��Ғ��i�  �x�m[��yMNN����i��E-,�k}}Mq7m_  �۶�y)�   @���   |�m���5���G�C�Ցp�ժ^z�mm1� :�������tS��5etiiQ�R�){  U�����ؘl�iʞ�W��Ғ���\D @�9��}��kI�    :	w   �s���|�����}��o�ǟhu$܁��^|�U*|�: t���~MLLjll\�i6e�R����E���(æ�	  �-L�����&&&��嚲gE*ֵ�0�b�ؔ= �.�q�����N:   �)(�   {\��}��~��������{���;�����/� �� �g����id��gZ[[���坦�	  ��zzz4>>���	9Ns��ߺ�peeYQ5eO  �;�u����N�9   �N@�   �d���A������{��S�e<��++˺t��* �J�411��ɩ&�bmnnieeYkk��   �a���ظ�����FZYY����j�ZR p�9������_'�   H�   {���f� ����̜�3�>G��������˗)<@�s���������Z^^���e)  �&K�3�����Ąl��%�q�Ba]���*��� ���0�ض����?N:   �$Z9   8�\��u����8�|n<55�g�;#�4�����t��u5rq �����Ȩ��g400Д=K��������(
��'   ~1�45<<���id����Ύ��紺���u  �a��8��yޟ%�   H
w   [�T�_�<��q|`c}||Bgϝ�iZ툆���w��;o' �%˲4>>����R�C�Ǒ��׵������&$  �������Ĥ��ƛrq��yZZZ����� hBB  ��0�T*�˵Z�GIg   �@�   ǒm�υa�b�6և�Gt��˶�vDC�|�u����' ��t:���)MLL6����յ�����y��߄�   8,�q5>>���)�Ӈ��1C-//innN�z�		 8�l�~����Ig   ڍ�;   ��u�}��8����f��z���$�u���X�_}E�|򳤣 ����ׯ��i��c2�ÿ�T,��0���5�q܄�   h>C��Ú��V.�k�~�
���~����&� @�3M��8���z�7�  p�Pp  ����d�����QeZ��ק����d\�6��PW^~Y��sIG�c����0������y���&�  @�d2=���h�7�p�#  �3Ms����;;;�Ig   څ�;   ���i�?��({��L&������׎\8��y�t�E���% ��i���ĉ����9�~�JE��KZZZTMH  ��X��|~LSS����=�~�jU�ZZZR�MH @w�,k#�S�JIg   ځ�;   �ײ�O�0�:ha*����%e��������B��t �j��jjjZ�r�P{�q���u-.�kkk�I	  �Ir��&'�522��~������0/��� �.cY��0��   t=
�   8L۶�����Z��?��FFFۑ�ժz�S��������	��c2M�P{�a���%��ϩV�5)!   :Y&�������eY֡���H++˚��U�ZmRB  ��m��A�s    �F�   ]϶�W� x�u�i���󚘘hG,�\.�~��߸
 ���ۧ����c2�ýE�y���5??� `�&  �qd۶���53sB�Tꐻ�*6t���U�}  nc���� �a�9   �V��  ��f�������0=��s��9юX8����^|�G�T*IG��30�Չ'5<<|�vvv������eEQԄt   8��T>����	���z�B����O���݄t  t۶�,�%�   @�Pp  @�r�|���F�>��i���o�:����_����z�Q ��d�Y��4��^,577�Ba�	�   Эx
 @�8��_����%�   h
�   �J���]��~����=��x�[��������K/�󼤣 @�щ'500p�}�8�����fU.���   �Aoo����466.�4���NI���Z[[mR:  �.�u����~�9   �f��  ���8���}�Y��C��G���Hh���.^|Q��' �����a�:uJ}}���)��,knn�o�   �������)MNN�q�C�U.�577����qܤ�  9��8����!�    @3Qp  @Wq]�W}���8�|�{��=:��3툅,..��˗�a�Q �H3S�|^'O�T&�s���ժ浴��(��g   4�eY���4==����=o�ժ�����Ң�(jRB  ��0"�u�B�^����   4w   t�q���8����NNM�̙s2�'mv���]�� p�eibbR��3J�R�ګX,j~~V��IL�  @�����MO���������j�������1  ��0�q��<��    �@�   ]!�N��y��Q��х</۶�_c��M]��2_% wɲ,��O�ĉ�r]�P{�E��ͪPXoR:   �q�lV33'5<<|�}|�������A�� ��LӬ�R�oV�Յ��    �E�   � g��Q8�k ���ˇ.��>���t��+���.X����iMO��X��뚝��R�Դ|   ��Љ'5<<r�}����ܜ��a�� ��,����$��  ��F�   G�cY���0�:ha&ӣ��/������5>��#�x�:�v �C�&��<yR�s���b�����O?U�RnZ>   �Yz{{53sB�����?��}_ss�ZXXPQt t?˲n�a�I��  ��E�   G�m�oA��A�R�����4�Ͷ#��G}��]O: )�ijll\�N�s�o!��H����y��J   ��N�5==���I��y��|Vt�WEML @�m�ZO'�   �[�  pdٶ��A<�:˲t���mG,|���Oo��F�1 ��0S���:u�\7u���a���%��ͪ^�71!   ���jzzFSSS2M���}Osss� ]϶��=���t   �nPp  ���8�����Zg��}�g�_�����[oQn�F����	�<yJ����7�y^   �pGSSӚ���m�w�O�^��ܜ��)� ���8���o'�   �S�  p�ض��A��F�>��Ӻ��{[	x�7��{�% :�a���t��)e2�����}-..h~~NA41!   �,�����N�8)�u�z�Z���ٛZ^^R�ML @gp���}��H:   p'(�  �Hq�����q|�s��<�~��툅����7��?M: t8C�����{Ul�l
咢(lb> �L�iʶm��%�4eY��cC�e�0ٶ��Y[    IDAT%ɐm����e���������6d�֗���{_~9bY�S����EQ�0��t�0��.e�{�C�q������� ����]E��߉�Xa�� �ݭ���̉C}�Ew @�2#v�x��'Ig   E�   GF:��P���<�c����}���O�#�ƍ׮룏>L: t0C�|^'O�ROO�]�R��t��M-//+�)38:Ǒm��7���c��|�fɲ�/��q�(���0P
�PA�+���,�ܚ�s?�� G�i���ɓ'�w_t/�˺y��Z[[kb:  �eFh��S���H:   �
�   8R��}���$���szrrJgΞ�a�t7I7n���>� � б��Gt��=����=|���ܜ���#��)�M)�reۻ�u�u�J���������9��<�.��{�'�����@��1�@������N��G�{��H_i������V�� �䘦YK�RT��٤� �?{w�����l��d�,�[w�i����H3�Όf�֌����q'���Ab �$@��͛8�� �'�vǎq� p�;�m�hf��Φ�H�n��fs��b�X˳�E�Z-���"k!Y�Phv���^P�S����   ��   8:L�\� s�����Wd�v3r�	(n�'������%�R��Q�V������e
�4�a�D��Ţ���"��"��'"�q(X��0��>(~���Z��\.�Z��R��R)�Z�@㙦���!����q��������Y��{uL @k�������Vg   ���   8�L˲f}�?j`*��+���X,քXx����'���nu 8s�ɤ������w�5\���ʲ��^�hW�w\�D�����b�G���(\G�}���R��\.�Z��R�<��\��@]X����!���ʶO^辻�����:88�c:  ���3�+��u
  �3��   8�l��S��~�q�hT��zS�tG3b�	(n�_�F566����������e-,ܗ�Q���,�R,S<W,W,{�g4��#�i�t�/�\.�Tz�g�\R�T� 5���}���BmnnjnnV�r���  h&۶��<��V�    ��w   �Y��������Y�����zzz�O@q; |�m;��аL�<��8۶?U�������bv��<�a����%�JeU*e�!)��z��a���5ݻ7'�u� ��p�����Z�   �<�  �L�D"�y�Z��G�3C_������HR�I(n�O������������Uݿ_�[�sB 珡X,�D"�D"�X{\�XT�q�M4�E��n��uxxH�e �$�q444���aY����=����}-//q� �\�m�?�<��:   �Y�  �̉D"�u�?�����^�M]��ڌXx���c�z{{59yI�X�D+A���5���S�Ja;�nL�R"XȞ|X������'A\t����=�~ ���� ���
�@��K
�y���?������g}��g�a���8˲>w�m[2�Ͼ�1dۖ$�4M��%�2e��uٶ��?-�z4����Z�%۶N\�y�A���Ç�E�҃�S�
��q42r���*���ߟ���*�G  ��0B�q�|�Z��Vg   G�;   ��q^�<�aZG���̳z���#C��'��ٻ�� -��եK�.+�L�h~Z[[������J��8k"�ȣ�O��'N�9�
�P���u]��'���y�c_�z�o�c_?x�h�m�eY�m=�ٶ-�q>��"U.W~��X,�u�V��`����ȩ
��������F�� �8�a��m��뺿hu   �c���4   θx<>\�Tf� 8��gttL_���6#��?�Sݝ�iu h����&'/)�ɜh~��:�W*��eYJ&SJ&�J�R�����U��u�uU�V������Կ��sG���8�D�:��=��__T��X,�X,���@�⁊��]��?�XL����r:�Խ�]��ͩPدo8  �4�R,�txx���,   �D�;   Ύ�i�KAt5���W_����#���A~�ӟhff��1 �e����'���w�5vww57wWuL�Ub���"�O����x�c�E��V��TʪT*�^�jE�ʧ����Ǌ�E"QE�^��(�)�\���J��c�:88P�\nu0 u�H$5>>~�{���m��ΨT*�1  �aYֺ��#�xs  ����   ��m�C��n5.�J�W_S,vd�w4�/���>��V�c @KD"��O���ąy������U>�W�t ���,%	%I��i%
��iu�	��Q�z�ZyX�^Q�\~��JYa�:*.۶�G��?�uD�hT�u>O;�}O��%U(tpP����ށs���K����N�O4?C��,���y6� �<۶�y���   P�  ���m�;���<j\4�+��T:�ьX����{��և�� Mg��4>>!�>Y�]�t�{��iss��� 4�m�J��J��J�;�J����A�\.�\.�\.�T*}���:"�D��(�)�)�+�)�?�:*�0[�w{/�P(�P�W�P��8Gz{�411y�{��p_��K
����  ��q�/�u�B�s   ��Q�  ���D"�u�Z���g�����o�/�kF,|�����n}�A�c @�uuu���)%��w]W��ZZZRR��U�a(�H��#�L&�;{B��#T���?^�^R�T��:.4۶+x�������Z�*��S>�X�~� ��8��P����'�DN�F�t��ٻ��ޮs:  �'���j�����  ��u���   �D"�J�Z���}�/k||�ё��������_�: 4U"�ХK��ݝ=�|�������������%�a(�J)�J���C�TZ�dR�qv?.u]W���_�Ǌ�Kt�>�eY������O^��:��a�b����{���b��F���,K��C�e�섧��]��ΨX,�9  �gF�8Ο�V���,   hOg��   .4�q~���ah5���׍g�mF,|����{����1 �il������NT�����V5?O�j�	��Ag�����S��L�lu�_�����cE쇏��]�mu<��pG�D�SE�DB�XLg�I��?x���U*�Z��<�����{���;ܻ7��z ��c�o��o���^��   ����Oj  p�%���R�t/��Qc'&/�w~��f���s�#��?ou h
�0��?���I9��:�nnn�޽9�΀��;{GGF�LF��]'��Q� P�\R�XT�\V�X��aQ�⡂�ou<�m��h4�d�A�{<W"�T*��e�7��\�����
������9�h�x<���	����h�繚�����2'6  ��4��dr�P(l�:   ��   h6ǲ�E��sG�������|&�k��۷?�{�h]]]�t銒�����y���j?_�d �bY�::��d:�����j��B�𰀽������CI��I$U:�V"�P2�|��Yy������W>����.ݠ�H�;49yI���'�xx��ٻ��ٮs2  Nβ�%���%�#   Ms6>y  @۰m����=wԸ�LF��rS�H���33���O�� �p�DB�.]Vww�D�Ţ���jgg��� <I$U&󠐽�#�t:���1���:<<��a�QA�����fY�����T�Lu{/�K������U,[	h�l�&'/=�S���-����d( ��a��;��}��9   �>Z��   m�q���_8j\4ի���T:݌X���{sz��s$6�Ͷm���ixxX�Q{�g�s5??���e~^d�R��2�·�;���R��b�@���\� �$��cJ�RJ&�R��b�x���Z�>,x�S>�����8Mh�0��?���I9�S��0������{�<�	 ���8�����9   �(p  @SD"��Y�V��q�i��/C}}�f��g,-.�?|�bM ��\.�K�.�qj/��Pkk��wo���@�$�Iuvv=|uʶ��)�K*
_�*
�}NeP˲�N��:�N���Z��u]���iooW{{�:<<liࢲmG����a��h�u]ݿ��Z ���8�_w]��:   .>
�  �p�h���j�����������ѥK�������w��=A��( �����|yJ�d�D�wvv4;;C�Pg�X\�LF�LF��YE�іe�V�*
:8xPо��/׭�,��Ͷm%�I�R�?;[zJ��V������]���U,[����ɔ._���ή�?88�ݻ����uN ���F��o���[�   �   h�X,6Y�VoAp�Y�7�yV�=�|3b�3�����?��H\H�HD�������h~�t�{��iss��ɀ��D��t���K]]�-�`�y����b�|>�r�Ԓ, �H$���{*�VGG��ȷ�Q�V��?(x���Q�\nI��f{t��e����___���,��  -c�f%�^.�JK��  ���w   4Rܲ�e���lM5<2��|��NtT3Ng{kKo���<�ku �3C�\N�.]>Qa��yZX����%N� N!����K������:q1�i�a�#����
�}
5��x\�t�����S�tK�;jooW{{{��ە�M� \�ahppH���m�����i~��VV��a �t�e���?"��B   4�C   h۶?�<�uuu雯�<�=�����~�U�t�p���i]�2�t���C����8!�0�J������;�t:����?,f�+��S>�g�
��4-��)utd��t*��m7����aQ���������E��	8����q�h���AA���*�� ���m�Ǟ���   ��(p  @C8��\���G����z�淔H$��)����7_�{)�Ŷm��O��@dooWw��U�xЀt���D��t*��*��i���j����}?�B�@�� څ�d2�T�A��L&�D"����kooO��[���V�Ri����.�J���+�d:O0���w9Y �t���C�u�j�s   ���   u�8����=j�eY��7_U6�mF,<�PЛo��R���( P7�\�.]�,ǩ��i�Tҽ{s���h@2��ie��0U**��?|�a >#�(��P&�QGGFi�ٴ��%mook{{K{{y�!�h Ǒ�����+��b5ϭV�������Z� �d���;����V�   ��B�;   �*�}�R������_���jtt���R�Po��]��VG��H�R�reJ��������E-,�WPx<M,SwwV]]����eYM�n��/hooW{{{*���~S� �eY��x�ݽ��K�tǉN�9	�����������`�511y���|~O33�|� h�0˲��y�[�   �   ��D"1X.�� �5��翨�7�iF,<�R���7^��~��Q ��,���Ą�NT�������YU����?�0��٩���J$M�n�:8(hooO������S� ufY�2�Nuvv���K�T�i��bQ;;����Q>��0�r]༉F����������a���Eݿ?�} �)L�,���b��Q"   �
�  P/�eYK����m||B/���fd�c\���o�����VG�S�f{t�ʔ��#�T����Cݽ;����$�7Ӵ��ե��^e�=�m�)�-�K���}�ڑ�yM�. ���;��խ��.���\��<���h{{[[[[�}~����٩+W��H$k�[�V477��uj �gY֊��c���  ��Q�  ���m���}�q�����+7Ot�2N��}�������F�� ����q]�<���������Eݿ_a4 p>9����z{����%�4~͏������vU�T~M ��9����.e2utd�R��������������1�ahppH�'�LmooW33�:<<l@:  >a��;��}��9   p�Q�  �Ss�t]��:j\<��׾�x<ьXx(������r�� �������1����0j/��������R�C�dR�l�zzz�Nw4�z�jE;;;�����U�_��$����K]]]���V$i�C���S�<��t��e�=5��@����� `�/ �q���\���[�   ��   8�q�5�u����Y��o|�Ue��&����}�Oton��1 ��2�N]�z�D�J���ޝ���v�牡t:�l�G��}J$��0Chgg[��[*
� ��b���٬��uvfN���rY��[�����ޞ�0l����.�����W��j�[*�4=}G{{�H ��H�_�V����9   p~Q�  �s�y��~��g#���W46>ބTx�/~�3ݹs��1 �Dl����%�<7-..ha�>�	ѶL�Tww���e�=r��׫T������Ύvww��~C� 8l�~��=���nE�ц^�u������֖vww��C�2MS��c�i־�d}}Mw�ޕ�H hw�ax�H��J�r��Y   p>Q�  ��J���A����o<���b32�1��K����V� ��f{t��ԉ
���v533����$�6�4��խ��^���Ȳ�]+C���?즻K�v ��Oww�d2'*�=� 𵻻���mnn*�\����u�򔺻�k�[�V533����$ �;�4�� �ćt   ��   8۶o{�w��q����^�ap��L��w�����1 �f�HD�/O������jEsssZ__k@2��z��=��m7���\.kwwG�����ّ�{� ��3MK�Lǣ�Db�Xî�y�����������!���^N�Ix{{[33wT�T� ��l�~��/�:   ���   P3۶���?wԸ���^����iF,<tonN��'�� 5���u��e�vm�7�0��ʲ�ݛ��ӵ��0Luww�����E���絵����m�J4] �\"�xT����Ѱ���ikkK�����Q��p�X����Q����0j;=��<���juu�A�  ��q���u���9   p�P�  ��8��﹮��5.��՛�R:�nF,<����w���<�p���q]�rU]]]5����433�b�؀d��b�:::��ۧ��\�6A���]mooi{{K�j�!� �7�q�ݝU6�UwwV�e5�:tvG;J&S�reJ�L��{{{�����F @]9���\����  ��w   [<�J�\�~�Ome�����k``�Y� i{{Ko���<�ku 8�0422���q�fm�]���ٻZ__oP:�l�tQ{�'Ґ븮���mmookgg��  Me��2�������)i��O�o�9^��.]�T�)Y��k~������� P�a�m���?mu   ��  �zMӼA���_��t��fd�C�|^o��]:�87R������褏����L�u�$ΆL&�\�_==���^*jk�A��|~_�K ��{��+���e�=�Ǐ��D\����66֕��r�,p��.]��\�������B�Ѐd �vc�f1�aI{��  ���w   �iYּ��#G�Ћ/}���P�t�׿�][ �d��FG�4::&è�c�r����;���iP:���ј���400ؠb�P����N�[* ΅X,�l6���>e2jģ�J��������T*�}}�,���jjjJ�h��yajiiQ���A�� څm�3��M�:   �>
�  p$۶��y�ͣ�uuu�Woʲ�fĂ�J��7�x]��t�p�e2�����D"Q��P������+���h�q��ۧ\.���L���P{{{��������  εH$������*��y��q��絾����y'�b�,Kcc�Q���K�����hoo�1�  m�q���_lu   �m�  �l���=��;G��F��y�[J�R͈I��������f�� �Sٶ�����yn�X���m���7 ��i���[�\N===2��W���kssC��� .$�q�����{www݋��0����ߧt��E��d45u�D��WVV477��c ��8���]��{��  ���w %��    IDAT  <Q<�\.� çV]���_���r�fEk{A����VVVZ ����[W�^S4�i^�ZZZ���=��pa��i�r�����q�:�NQ; �}5����<mooi}}M��t���`���G411Q��r��;wn�� pb�a�m���?ou   �M�  �I:M�\
� y�����4u�Z32�w�����Ͷ: <�iZ��Ȉj��a?�;w���ؘp@E�1���i``P�x�Ϋ?^Ծ�j�R�� 8�Ѩzzz��ۧL&S��+��666����R�T���fK&���������箮�hv�.�� 'b�f!�AI��  ���w   |.۶�x�7uԸ��	��җ�	���/t��[�� O�ёѵk�k.�_���ZZZT�J4�eY���S��::�_X�����Ɔ��6U�P� ��D�Q�������DŻG���Z[[����8��ҥ˲,����rI�o�V>�נl ��̶��<��R�s   ���   ��q���xԸ��.���MY�݌X�t��~��?mu �\�ij||B��#2��>r�������*�r�����ѡ��A����\t����;�oP� �	�b����J��[����66ֵ���Ba��k���45uU]]�5�������YAАl ���q���u���9   p�P�  �Oq篺��?5.��׾�d*ՌX�������}�8���]�v]�D��y��innV��+J4�m��������Ru�/�T*���J�ú� @;���}``��S��rxx���U����uݺ�4Koo��\���85�+��s�#
�% \T�H�/U����   8;(p  �#�H�Y�u���-G��W������moo�7ߔ�{�� �b���G411Ys������LS��s)�Nk``P�\N�Y�n��i{{K��k��ݭۺ  ���i�r�����\��4Ah{{K��+�Nǹ�D49yI�\M��0��Ң�ݻ�0��; �x��"��3�Je��Y   p6P�  ���M�\� s��/���z�Z32A�A���_��*�J�� ���R)]�vC�d��y�JE�ӷ���Ӡd@cD"�r�u�������������M�_�� �񘦩��n�r9����0̺�]*��ʲ�{{�;�l����*��4�P(�Ν�T,� pј�����j��   ��(p  �$ɶ�_x��ţƍ���/�����x�;<p�|ҵ}����MOO���ڎ��PWW����[�IOS(�������.�n 8+l�Voo�r�~e2G�8��7����hkkSa�mm��l����%�4/C-,�����|� �Ŷ��{���V�   @�Q�   9��?����5.��ԫ7_�m�͈��<�՛o��Q� ΔD"�k׮)��i��V5==����%�+�i``@���F�u[�\.i}}]��k*�Ju[  4F"�P__N�\�b�X�֭T*Z[[��;Ε��>]�2%�qj�����;w>���a�� .�H$���j�o�:   Z�w  �6�F��j����a��{C�qt��k��_�2<Y��������VG������2M����������ҵg_WW�����ԭ[��y���������|]�  ͗�t*��W__�,�>���0����VV����s�q"���ROOoM� ���=-..J��; ������7����Z�   �C�;  @K&��R�t?�#ے~�wO##�͈I��cݛ�mu �$�b1]�z]���5��<Oss�Z]]iP2�>,�R__NCC�J&�u[�P(huuE��}�n� ��2MS�l����U�uK��VWW���"���.���}����m���=���Ν�8� �T�i�� ����,   h
�  ژeY��5���z��/5#$���_��?hu �$�r��reJ�U[����MO�V�RiP2����400(ۮO֏��///�X<�˚  ��J$��P�'R�5}���ƺ���T,�&��HDSSה�fk����fg� �T�m��<�z�s   �5(p  hS�m���y�q}��^~��2n�anvV��?nu �mۺreJ}}�������Y���,3��f544\ǎ��vw�������AP�u �ya����������[��Q����������0�&Po��t�r��7774=}�  O�8������   h>��   ڐ�8�u�xԸX,�׾�m���f�j{����oQ��:;�t��uE�њ�����Ν۪T�J���D��߯��!�b���Y�V�������˥��	  οh4���\��;�Z__����$�L��b�z��:;k�DZ.�u��G���� p�E"��Z�����  ���  ��D�ѩj�z+ç�T2MS/����6+Z[������U�Zmu m�0���ktt����Ah~��%�UgK:�����r�~��y���0��ޞVWW�
  �`���S�u��������������:d��$���0��Ң�ݛ�� �k�p���T�\�ou   4�   ��6Ms5������o����fdj{�rI��;*������b1]�~C������u��m�J�J��0L�r}Q*��˚�RIkk�Z[[eC  �Y$Q�����vR��AAKKK���PrΎx<��W�)��i����n߾�R�ӑ  �fY֚��C���  h�  �۶��<�w�7:6�/��a�����[oh{k��Q ��\�_W�L��a���KK�t�Ùaێ544�H$r���0����VV��
  ꦫ�[��C�f�u��^�V������ey�W����������O�t���{������z� �#۶���y�B�s   �9(p  h�m�g����G�����͛ߒ�8͈���0�����[@��m[SSW���WӼB��۷o���8b�������?P�F�'�<O��kZZZT�\�CB  �_�D588���!9u���}ml�kii�{u��TJ׮�P2��i����ff���~�� �#�q�C�u��V�   @�Q�  ��y���a���?�q���o)��Ѭhm�?���ܹ�� �TGG��_��X,^Ӽ��%���*9��N�544���\]��
���h}}MA��8  h�0��ӣ��Auuu�a�P��;Z^^��	�ij||B###���t�\��۷��� p��ض����:   �w  ��/a��Z���җ5>>ьLmo��]��'�:�6d����5::VSAp�Z՝;igg����0��f522�L&s�Ղ �������(�  -�N�500�\.'�<��4�BA��K��XW�uH�\WW��]��H$r�9aja��ߟ�{  I2Ms/���j��   �q(p  ��l����y�qԸ+W���o�V3"����}����C9 M��t�ڍ������4=}[��6(p4˲�ח�����ĩ׫T*Z[[�����  �̱m[�\���G��N�^�\��ʲVWW�y^'�8��^��l6[Ӽ���>��#�˥% �'�m��[�   �C�;  ��D��j�����ݝ�+��Z��`x���]���wy���z{�45uU�m{N������R�O�D488���!ٶs��vww������M6� �s�PWW���Fj.�<��immM���T*u������._�\�瑞�iffZ�L 8/l��O=���Z�   �A�;  ��8΋���(ç��E"�|��J�Rֶ͊J��^������Q �˲555���\M���G�3-�L&522���>�y��|����VV�U*��  �O�xBCCC���e���	�@Z\\P�X�SB�6�dJׯ�P2��i��ڪ�ޝ���J 8�l�~�u��Z�   �G�;  ��7Ms=��Q������fdjk���7_���v�� h#�TJ7n<�x<^Ӽ��%���*�%�,�JixxD�\N���Z�juuEKK���  .˲��?����b�S�������y����!P�459yICC�5�;<<ԭ[�A ڜi�{A�$U[�   �E�;  �d��O=�{�q׮�����fDj{?���p�~�c h#�\����j:�Z��Ν���a3�/��hddL�l��khiiQ�
ð�   �"C�lV��c���8�j�|^����ުC6�6]]ݺv�"�ȱ�A��wg�����d ��ζ��y��r�s   �����   �B$�ۮ��ţ�e{z��K_�a�������;3�� ڄeY�v����e������W�����u]]]�~����&�H$N����fg�jv���E�� ��W*jmmU{{��,K�D�ğ��b1������-�uU*�9-�d�rI���J$��~_`�����q�� �T�m�� �a��   �~�f  �@�y���a����H$�׾�g�L&��m-,�׏~��V� �&��n�x����AhnnV��KL|փn�cccJ�O�m4mnnhaaA���:�  8��񸆆�500P�iN��X,jqq�Sq�tCCÚ��$�<�����Cݺ���E� @;2#�m��u�ku   ��   G�4�� �Od�����k``�Y������z�A��( �@.ׯ�����X�Ţ>�����4�a��/��ѱSwkw]Wkk�ZZZR�Z�SB  ���q��hxxX�H�Tk��%---iuu��8�4�dRׯ�P2�:���5=}G�L 8�L��� '���,   8=
�  .۶�y�o5�g��/|�fDjk�bQ���T.�[�g��._����@M�VWWt��]�ߠd�'�T__������O�V�T���VWW��  8�i��������O�+��ZZZ��Mc��&'/ihh��y��k����� �!۶��<���  �ӣ�  ��D"�_�V��Q��r9���7e�6��z���h?�ou \2�ԍ���	�u]ݾ��vv��x��,ixxD�H�Tk���iiiA��;���  h���n�����T+U�U---jeeY�O1���WW�^�m�Ǟspp�[�>P�Tj`2 �Yd����<��:   N��&  �s�q�/z���0ͧ��F��ַ��SwM�Ӆa�w��c�,/�:
�.��ו+S�,��s
�}ݺ�!�K��,��������e�Ω�������}����)  @{�����蘲ٞS��y����D�;.��ƍg���q�9��kz��666� p��8��j�z��Y   pr�  �o�eY��w5�k_Y�����~���jf�N�c ��NzD���fgg�A��
���4::vʎ��wt��=
���  �'�ɤFFF�ח;�i��jeeY����}��	�O3C��i�������(x? �²�M���%��  ����  ��m�m��~Ըk�o�_�R��{ssz��?iu X"�Ѝ�(�L{��y�������&C�3S����8Ua{���X���}�1!   �$�ixxD�2ͧ�T��jqqA��K��zzzt��uٶ}�9ݺ��J�R� �۶����l�s   �d(p  8����]���G�����Wo��%�������z�� ���WSS�jz�_(<x�_.� ��qa��ظ����	�@��k���*�r  ยјFFF400 ӴN���V���H�;*��ƍg�Nw{��{�s�677� p�8�󯺮���  ��Q�  p�b��J�2��S�#��^{��J�����+�z���r��< �g��&'/ihh��y��+���QRP��3C}}9���+��x��������U��:&  �I9����a״���*�����B�;��� ������b����ÕVg  @m(p  8˲}�:j�K_����ƛ�}���7���vvvZ�����3_P���J���Ν����l`2�/C������T<~��v�u������%y�[�|   �˲��?���1E"��S��u��}���*�:&���ij�,��'������� ڀeY��O�:   js��  ��m�S��_<j��+Wt��3͈��~�'?���Z�c ��:;;��s��TD|pP����R���&C{2��ۧg�}V��Cr�D��nUKK���[��١�'  ���
�}����Z�*�L����m��f{���+�H�vV,�������coƈFc���W�P�TF ���0�tg0���,   8>:�  �#�H��V�����q�L�n������v|�+}��[�400�+W�d�۾����wg(F�=��>>>�D"q�U*��t��{  �|2M�QG�h4z�u5?O�������1MS���444|�9a�޽9-..40 ���#�ȟ�T*��,   8
�  Ώ�i��A<�	�mۺ�ڷ�ёiV����������PW�ijj�r��c��}_�ӷ�����dhG��YMNN*�L�x�j�����Z]]��  ��0MS�;v���S,u�ެ�����r���\�ZS󏍍uݹsGA�70 ��L�,A�/i��Y   p4
�  �	۶�=ϻrԸ�y�%MLL6#R�������ߑ뺭�����z�/(�L{����n��@�R����n��MNN�����k�����-//S   pA���\�_���*t���knnN��^ӡ�%	ݸ�l��?��W*��L h%۶�y���  ���:   Z�q����o5nl|\_���͈Զ*���z�t����n=���Ŏ=g}}M~��\���dh'�XL�/_ѕ+S���'Z��\-..�֭[����  �,C����j��T*]S��E�1��(����A����u����H$�t:}�9�HD�\�
|� T�H$�}����  ����;  ��8�o{���0�z�J��ڷ���iV�����~�Mm���:
�dttL:�[� �u��ml���8�FFF544,�4O����ZYY���}y�W�   8,�����FG�d�����Pkk�����j�ͼ����]�<u��;ajnnVKK�N h�0�q�X�V��,   x2
�  �6�4�� :�6�0}����iV�����T��wZ�aY��^�����cϩT����T(�������1Y��
�(l  �gգН�L�[*��3�<[��i���-��� �
�em�����:   >_��  �il�����7���s�kl|�	�����y��hu D<�s�}Q��Oݿ�){{{z���T*����0�g�����um�}_��+�u�Cmmm)x  ��0��~^���
�@�t��{N�4��d400(I:8((�F�E��V���XW*�V<?֜d2���vww�h L�	�qnA�O[�   ��w  �3�q���y��8j\oo�~�w^�ap8O�����w��0�x��e�Y}����5nqqAw�|D�8�Zoo��y����e���PZ[[Շ~���M�'  �DAhooO�����t:%è��ݲ,uuu+��W:88hDT�� ����h�qD"���tpp�r�� p�A�L$���g��b#K�41�g���sg&���Yj��-�$�ZR�Jj�g�i4fు_�¾�Kc�r`����� 6lx؞�ѪE*Ui�Ekfrߒ�=�q�,�`f�RU"O0�D��d~��� V�����a�w:}�����������T*��i��թ��o��m�|�vE�9�z��.�� ��Z`l�&&&`��a���@2y�l0��B�0&&&�]k�eY8==�ӧO�i��#"r� �$	�(B%H���{Q I2A�,K �g���LY�?uc�,˟��eY��	H��OL �x�i0M�qQ�� ���z�����&RUw�chh�ڃ�������e[��zM� fgg!��6�Z��������p2""j'Q�i��"""�.�w"""�.$����W�}�K��Ν��ԓ,�~��D��Q�膓$	ss����T�U��>F�\v0�v>���D�׾F2����*�J�]M�$ȲY�!I2dYz��'����o��_4��V�i�4M��w,�    IDAT4��:t݀�7^�i���0�������</�ݛ@<n�����d������%z%~����M���N������c(�m!��t]�l�s����NDDD�eTU�ך���Uu��S����Q;"��_������t"��^�����xm�I����Xc�]�,+���ȵ�c
���"�ϵ8�*Q!�
\.��zќ�r���*dYy�w.����)��z�iB�u��uh���A��ס������'&�]W Ї��	�B�k^�B"����.��٨w(����E�����2VW�Z�:�����IU��i�_v:�܉������(��u��-˺�y�?�[�z���+Z�y�������v:�p�p��e��������`�5O�޽	(�|�P�T�����y���m�(ꋦt��UU�v�_�\Q(�z�7�]�Ƴ/���^���Ҵ��k�,��Q���Ø������z]�qp���G0M��P�A��{�c{��7����\.�`2""jALEQ�5M[�t""""��O������,Iҹa��E_�ƛ�F����s��,����y�0����aLO��n�3�H��'��*crr>��Z���:�>����)���3³�u����n�E��&���N����]���j/5�?�Q����qLLL��v_�
�jO�p�&]_<ޏ��9H�d�޲,��l�����dDD��$%�'�u6�u	Y������W�}�3�ٹ�vD�I�����A�T�t"��A���FFFm��V+X]]A�\v0�V���S���f��qp𔍆D=HE���n��n���^��v��u躎j��Z��Z����j��Z����A1<<���{M���q�l���|}E���z�����k{���	����Q���P��5���DDDD�w"""�����?�4����nppo|�O��'Y���>���NG!�J�,.."��0����ill�A�yj5G�eܹs�����'[����3<y����@B"��n׳������7�+���D��4͏5��n|����n���uGFF�uR�eY8;;œ'{h4$��L�d���#��^��d������DD�����v�^��9����z܉���:/(��i������*�z�;MM��<|�k���u:�P�KK����><<���8���#``` ���P��-$�I���V��<u� ��z=�z}p����|�z}��N���i(�˨ժ(�˨T�/����p�\�{w��C��?������qrr���Դ��;����ݏԫ�
?~�j��l0""r�(��4��8"""�b�;Q�ɲ�+]�?sU���:�ܹێH=���?��G��AD7T8���dY�U��:66֐N�NF�M8���4|>ߵ�g2���\.�8������z_��x�p�/�/۳,˂a0M�i�0L��	�0���˲�����瞯�]����À �:i�Ӟ#����A�$IE�(B�$�Y� P�Ś��I���R)�R�|쫌Z���V����cbb�H�Z���2vw���f[��n�X,���yۏ��F������NFDDN�e�������DDDD���DDDD�(��h4�����ݛ�����'��E���;<����ehh��3��	V�U��<B�nd�����{������Z��ɓ=$��-NFDN�e>�>�~����^H���T7��FC�a�/��u�ٟ��z�����0L�����=o��e�ŗ$}�{����Okȿ�,�D�RE�RF�TB�\B�TF�^�t4"j«n��f����F��d������}�
-����&���NFDDNR�_6���DDDD���DDDD��x��j�]˲.�P��|x���@Q�vE�)�a���{����i� �޽	��ݱ�&��cu�17Ԑm�$���q���B�o@�uO������Sk�������z�����^�q����	M��^מ5�7�i��������hh��j��y�"CUU���,CQ����r]|��CG�TF�RF�\F�TD�Tzi�?uA022��w�m���q�e���O����u�MQ,,,!
�^s||��� |NCDt	���z�w��2w,u ܉���:D��'�a�_V#��'_G�@�R����ۿ��'{��AD7�$I��_D4������ۛl�#ۢ����mO	|��D"���]h���lDt=�,l�~�>��(u:�+i44�����u��5��4��F�Mk��]��$=o�W��.�\��RU�n7TU�}�M7�,�j�ٔ���2��j5N{'�&��`||��#׺�Ѵ:����H�g��E�ӳ��&�Icmm�'N�!"��dY^�u}��9����z��}������SU�_k��W��/,������'mom◿�E�c���x���l{��eYx�d��'�����`jj�����e����R���dD�Q���������b:�M�ij�ڋ��Z��b��󟙦���u�����K��u��~���u�Ӛ������⳯7�u�׋�ɩWz�����J���dt[���bjj
v?j/��XYyčRDD7����JӴ��t"""�^s��=&"""�TU��h4~mY֥纇�a|�ͷn����"�N����8DԔ`0���e(�b��0���!�N9��nA1::���{�z����x�(�:Ax�^���gM�B�?��,�z�j�Z�j�����J��F�Q�,��������v����q���t:�-���X,�T�hz/�h4��Eԓ��&'���4�aYNN�����p �6�H�$�V}�����
����Ɉ���A0UU]��뛝�BDDD�K��NDDD�^�$Ig�a�/+�$	�|�-�B�v��)�Z��'sQS�033c�Y�V�be�1�����6�����tg�0ptt����ܸE�ϛ��>���]���h4P�T>��^�V9}���$�/�/�/��z/���7���K��K�"f��D�`|�d�^����jU��l#�N;��n�Ϗ���g�KW3M[[�ܔLDtI�tb�H�s���}�����R��Ɵ]U���fff���X��~�!��N;��nA011���1�k��VWW8�����.LLL```�Z��3���A��A�$�����/�`0�`��l�$�v�4�r�Z�r�J��dv��DD�\.�|>x�^x<x�>��~H���x�`Y��
�����j�Z�c�j�����q�@��84�Ncgg���ҕTU���2���l�98x�'O�LEDDNP�j4�e�s�
6�����z�^��wU�����ڟ�#ROz��7X[[�t"�!DQ���<��~�k������$m���ɒ��M\��X,`gg�B��tD�MUU}�����/�U��M�|��^��^4����&'D��>�n��Y���$�n�i����<J�"
�,��t,�[���cjj�`�$����C��DWE33�Mm\N&���X���"��v�_�V�?�t"""�^�w"""��p���2M�Y���x��߁��mW��rrr���N� �B�,--#�^���>���8��n�P(���x����jZ��;8??w Q/���_4����N�z�B�ZE�TB�\~�g��d��I�e�|~��~�|��bwL|7�|��Ŕ�b� ���V���199�����J����-�rY��m26v��|�����c��FDt����1M� ��9��DDDDm ��{���yU���:�ܹێH=�R��w��z���(Dt��,/߇�koÑa��XC*�r8�d��bbb���~�Y����c<y���;���7� �?�P(�P(�`0I�;���h`�m3{�ى'����Nӻ�+6�X��R��|>�\.�|>]�s �W!��ܹ�;w�\�t�t:���M��D���㘛�����R)���G��HDt�(��W�F��;������c�;��TU�����?WՍ����/��z�i�����T2��(Dt}X^^�������:VV�T*:��n.###�Yn��6��c{{�rɁlD�� �߇P(���=t��[�b*{�EC{�TF�Ά&�n�������b[�Ὀ\.�l6�|>�M0D����0==�`0��Z]ױ��''ǰ,ˁtt��~,-ݷ}b��ix���W "�A\.כ�z�{��ADDDt��������YnQS�i�.+�x<x���\�d�گ~�Klmnt:� �X���'�
��>��i'�����aff}}}M������q||��3Dv����a��a�Ba(�ұ,���X,�T*�X,�Pȣ�ht,]� �z�������\k
t+<���e��f�5���BtSbbb�jos�ǕJ%lnn�!�~/Uuaii	���ׂ�a`mm�L��dDD�
�(Mӌ��|""""��������A�,���W�}�o`xx��z���~��v:� CCC���� �{��L�ccc��D��A������]k�k"q���6�٠�.�A��aD"�\���u�r�R�|�|���n9A�����D p����zщ�^L�D>�G�pq����aY|�JtY�1>~��#�_>gY��������S�����9��ت�,��[8==q8��,������I�s�Vlp'"""r����iڿ��nrr
��?jG��S*��޻�es ]i|����]xx���]�э�����,|�Kp�T�R	��[(�$#�$Iz6�=�H$
����i�P(�X,<�*�V��=uY��5��!��������t]G.�C&�F6��}��~?��g�u�R�Z���&r����6�{DD�����PӴ���DDDD�܉�����E��4M�eE>�o��(�Ү\=�4|�����f:���� ����45jQ�0>>��ѱ��?꺎��'899�eY%$���n��(�����NFx���X,"�ϡPȣX,rR+�����`0�lڻ��x�V�"��"��hx�}ѧ000��ɩk�Wwzz���]��@6��=5���[[|}HD��DQ,����DDDD-�w""""Ȳ�S]׿xY� ��׾��{M�Ԝ���ﰻ���D��$I����ርz�0����t:�p2��"���g�5I:�<���64Ms ��$IB�0��("�\��Ni�ժ������(�(��m�}"��$IB__������ �R�n�4M��yd���iT*��#�8YV0>>���4�Q��i���B*�t&�h�X������,VWW�i����ɲ����ou:�m�w"""�S�?o4��Uu��s��|��z��ӧ���~��D��TՅ��������5M���#�E���M#�2&&&144���j����m�6B���C$E8A(� �gJ�eY(�J(.�s�,�F[n���� ��z�5�
�ں���t�l6�L&�0�v�D�,azz>�����9����hp+�,����2E�U_.����#��u��ѫPU�k��u:�m�w"""���E��4MץE}}��[߆$�oB[�(�x��w��lDD����ay�\�K�_�T*x��!j5�2K/�����4Eij�i������C7O=M%D"aD�1D"Q���&�We�&
�r�,r�,
�",�l�m���x
����z���J��N��PI=O���a||���vww�H�9��n*�ۃ������ڪ��jx��!*���Ɉ��DQ����㑈���Z��DDDD-$���u]��e5� ��|�h�]�z�a����!��v:
u�p8���%Ȳl��P�ce�1'��KTՅ���b�?���9lmm�1�z��(�D��F��D�m���|B{.�}1��Ӊ��q�=��/�d��v�U���N��N�����r�D���vcff�p�鵹\[[�V�$��JQ,..#ڪ�u++����NFDD�%��G����9����n6����(���h��W�-..a���vD�9����cgg��1��Kbvv�`�p*����L�S}鷆��199�tS��������c ��N���v#�!�!
پ�>�J�|�l�l����-#���/���=b{竨�j�f3H���d�<��zR<ޏ��k��d`��8�KDQ���A(�ibss���'#"��RU��5M��N� """���NDDD�}�(���麬(
��o�Qە�g�?�q�cQ��s�.�ݛ�]tt���]����z����C_���z�L&���M�HFԍ��������z��J��l6�\.�\.ǆv"�)� ����P�P}}A��wh4�d�H�R�f3<�z������F<����B����u��D/����i��\aawwGG���""��E�j�f@��Y����n:6���,����]V#���[�D�?ʘ.W����;�e� }���I��ݱ]�������Msݩ횦agg�dҡdD�CD��a�b��UUu��CG6�E&�A&�A�^s����nI�
��DG��x�=�4�MvO!�J���ks��h�ӳp�.�w�	�ib�	���KFFF155��`oo��PDDt-�,_��ov:�M�w"""�W����i��~U���2���#RO1M?��{H�R��BD]F���bpp�V�i���XG2ɣ�������B�p�k�3����h8���;<����� ��8z{�Z�t�t
�\�e:z{DD����A8F8F$mz�^s,��$��H&Ϲ�n=I�q��=����ُ]�<666P�r�;]��㘛[�}
���1�����爈�����HӴ���DDDD7܉���^�OŤi���C�Bx�[o;~Dx/�ͯ����N� �.#�"����m��z+++��s'��b``��3M7��jUlmm"��:����^nj87��0�r9��)d2i��u�n���W���`0�p8�P(�@ ��mY��B���������V�������mj��i�`�2@(���dY�U�J%������O"�n"�b�4� 9GDDDtMlp'"""z�,�H��/_V#����D��g�����}��D�e$I����ር�Z��Ǐ�R��<TU���,��XS�,����1�<كa�#�A
�������^,�ɤ��dP,`Yl�""r���A$A$E(rl��eY�f�H&ϑJ%��#�C�I� `tt��݃ 47�"��bss�:{���|X^���m�>��bu�1_�uY��Z��?�t"""����DDDDפ��i��WW�-..a���vD�)�Z��ר�����,+X^����>[��b++��i�&I@<ޏ���rsͻ�r	���(%#���Ť�x���̤��O�M����ND�Aϧ�G�1�bq�\.Gn����	4Gn��S|>fg��{]��a�������C��&QU�����m��<~����DD]��r}�^����DDDD7܉�����-�b�4�K����[o����^eY>��H$�:���������l	�ɤ����	gEQ133�X,��:�4qxx��O�²x<��`�����Pg��u]G&�F*�B&���0QW��ׇX,�h4f�9v�L�D6�y��)���Earr���3���6�� �2�
�m՗�%<z��������(�E�4� ������Ilp'"""�Y������/�����F��g��<���G��AD]���������>?O`cc�e9���]<ޏ��(JsS��66�Q�VJF�>n��x?�����x��Z��l6�t:�L&�M!DD7���A4E4C(� ���%�4�N��H$�ɤ�\�n�ǃ��y����5��l���ܡdtS��������6d�j5<z�T�U���]�,�ߺ�����ADDDtӰ������I.������xU���"�?x��zJ2y�|�}~�MD/,/?�ݠ|rr���m ��e�,cbbCC�M��,O���>��F�e�x?�n���R)#�N#�N!��;rDD�~�� �"�"�:rj��iH&ϑL��1�n���aLMMA���%�Lb{����    IDAT{����2A0==���![������(�J'#""��n�7j����ADDDt��������9�(�i�4����x뭷��Њ.�i�}绨Tʝ�BD]"
aii�$۪?<<��ޮé��E"�����r5��\.ccc�Mtc���h4���AD"QG����y$��H�R��k-�>uI�G����iv/�KH$H$дz˯O�.^�ss���Z�hh���B*�t(���c�V�u��<�&!"�.!�b�4�( ��Y����n
6�5A���O��?��F|��B4mW����O�v:u�h4���%��h�~wwGG���n&I���18ho��s��N7] ��� ��l�vьJ��d2�D��j���'"��A���X܁fw�|����0���#�ܹ��w�B콖}.�8���6Cw(�ccw011i��4��� ��8�����P��h4���9����n
6����x^��j?�,���P�x��3��3vww����N� �.100���y[Ӈ-����&��Nې��U ���"<OS�*�266�Q,JF��ǋ����v����B��9��$'��'���h4�x��h��'���T*�D"�\.�M�t��|>��-�����O��j��X�T�7<<���i���߲L���#�<w>]JK���7�_t:�M�w""""{Q�ώ���>����9������;�uN�""`ddSSS���4M����(�722����&'$Z8>>���.L�t,Q+���h4���a���_��ډ��:���iu$	���V�+�9A����ݛ��y�9�0E ��1?�`�T;˲�����ӓ6$#"��H�tj�p�s�lp'"""�AQ��h4��e5� �O�������L����t��Q��4s�aX]}�l6�p*�V.�ss�BM������|>�P2���z}���Ei��Ԟ@�Zi鵉���8��n!������T
��M�t3}������mj]�P���7��p8���e��������u8]EU��NӴ��t"""�n�w"""�+��:�h4V-˺�����4>��Ϸ+V��ͯ����N� ��0==���[ՍF�=D�Tt8u�X,���٦�}OOO����0JF��$���CC�-�v�Z��y��ډ��Q�$#�a``�p��Ȫ��pvv���ST*ܠE�OE������XS��C�������n�����}Ȳl��M�DD�'��r�&k��~��u36�]A����aܹ������o�)TUmW��pvv�~�!�[&�yfgg188d��^��ѣ�ld�Q�(bbb##�M���j���@.ǉ���� �����?�ҩ���#�N!�8��DD�v��B<����~K�],qzz���71R���bnn���u��9��6��Cɨ��|>,/?���Uzz���- |ϕ��SdY^�u}��9�����܉���.����i�_^U��/#��5�����:�}�95���	����9ڪ�T*x��7���'�n0?� ����:6�P��e�x?FFF���ϲLd2Y$��H&�0M6�Q��|>b``���C���9NOOP,�'�^�(abb�Z�v76֐��JF���v����lo�8==���&��ND�9���7�F��t"""�n�w"""�����T*�#˲.=����q|�_jW�������G��ADt��>���[��b�?D��p8u���QLNNBD�k�677�N�LFt}�P��#��bM�n_�P�#�H������L""�N�  �``` �X�غ�K8՝n�p8�����6zX�����x�t�'"� UU�����I��	ll��w���CAhX�5 ��,DDDD݈�DDDD��,�u]�Y�������S���v��	�[���/��D�A� baa�X�V}.����c'p�UU1;;�H$�Ժl6���uN���#�"��~����tZ{�^{1��'��M#�"���D ��x��T���#���\������N4���B!���5�j5��Q��eKK�m�'��X__c�;Q�Ȳ�S]�_�t"""�n�w"""�O�(�?o4����?��1>~��zF���{��	jD=좹}�X�V}:����*L�t8u�X,���9(�b{������Q��M�^/��G000Y�� !��@2y���S
��\�����\.188��Ӳ�f�#�N����cjj���t]�����&�n$���Dl�'�I����ɝ��CTU������N� """�6lp'"""�$�(�)�4/�>44����ve�	�i���{�Oc$�U�(bqq������677�!l�E	SSSnj]�R���J��CɈ�% add�驜�)�H$ΐH$�덖]�����c``�������u�������G�{�|~��/���5����;;�&�cA����q{'�R�,�����MŊi�Q <z�����c��NDDD�;dY����v�˲�����~�b�������N� �E	KKK��5����bss���[�^/��5��H�a{{�M�dY��� FG��v_���6]בL�����R�%�$""�)dYF<ޏ�ᑖ�Wc�&�����x
uQ111���Ѧ�U*����\���^"fg�000h�>�Icuu�'�u�,��A����DDDD݄�DDDD�r��Y��߿���gf��g��I|���8���GI����e�Ba[���'�����{K� fff!I��s꺎��M���;���'���E��� �H�4��������m�@S�/����36~RW�#�������ט����]9���� ����࠽&�\.���G�ND�~�,�_�u�o:�����[�������QS�i^::8����x���R��h4���E��F�z�Es�}�B![�''����r8u��N)����XG�^w(��A@<ޏ��Q}-���i8;;���)��jK�IDDt�H������1���pzz���#h�֒k]������C$mjO��M��3�U�����1�܉��M���a�v$��֌� """�E�7�a�~Y� ��W߀��iW������=����AD �2���`�V���vwwNE����������l��,O���	]�LG��I����,,,`pp.���h!���ɓ]loo!���������e�T*����T
�e���B�k_S�$�!������V���h�05�}�i��<]�
�m���������s���!�L������?n��`�d��S+���Ų,���n�0>�t"""�n���DDDD �n��z��cY֥�r.,.�����������1��.��؞�xxx���]�SQ7��☝��,˶��j5����P�;����SU��#m�w���u�����P�qZ;ѫE�h��c��<����8<<@:�j�������a~~>����4������S�Q������蘭�b��G�B׹���]A0<ϝJ�r��,DDDD��w"""" �,o�>sY�������Ӗ4*хZ��w��k�j�NG!�6S����އ�ln�-�(bbb##�M�K$ΰ���cԩ#�~?FG���?`{z�eJ�"NNN�H$`���&""j�@ ���a��T��������H��49���U^Gmmm�9g���w�mՖJM��OD�>�,�J���v:Q�I�@DDD�i���K]����������lG�����l��1���TUŃ���ܾ����ONE����`y�b���5��cccOaY���~��p8���LNN����Rs�e�H��������J�"�����i��4��N�h4��z_i�����Fc�,�(��lt���,�L�r	�H����ߏh4�\.�I�="���4M�Ñ+kUՅp8�T*��4"�61MsHQ�'�i>�t"""�N�w"""�u^QӦi�/+�;>�/|�K�����6��_���1���TU�������٪�����ѡé�[�b1���7�XT*�����j��`2�����x�w�܅��}��i��D���G���-HHDDD��F122�p8��W3M��9��R�� �}.�M�0[[�8?O8������LLLڪ�T*x����4��TDD �(VLӌ �EDDDԳ8�����z�,���1sY�����W�x�)^��b�����'�,N�!�%���k����f���-9���� �����Ԍ�)� �H�auu�?`��Pw�����"�(�+]/��boo�ۛ�f30�EI����:��
�3�RI ���k����	� �ߏ���|~��und��1��DQD0h���bg��L�'	��B!o{���(�F�H&�0M�n!"r�eY�,��i�U��u
'�Q�r��_��j]U����1&&�M���Y����}�өNG!�6R����^{�۷��prr�p*�.���,H]��rattCCÐ�W�aƋi��JDD��$I��� FFF����-�\O��f[�����EW����3`^(��x���h4�"""A,Y���h4���Y����:��DDDԳDQL����&��׿��vE�	��+x��a�cQ)��>����v˲�������6$�N�Fc����,۟�].������`j��������[��4��'8>>b3э# add�h���V*�ptt�D"�S��y������躎��$�I�Q������J%<|��:_�9M��S�0�;������^m���(��h��Ո���~����6���r�,��o~�#��z�,˸�5���+k-������6$�N����Y����&�3���@�4�>���S���C__�p��r	��O����l6�4[�����ڥV���<�t:I������AUU�bq��q��J���D/�u��dYF__��5�("���B&�q8!uZ�TD�^G,�UM"� �<��""�Y�PUU2��Ng!"""j7Np'""����z����eY�v�-.-cy�~�b�z�i����E.��t"j�������ܲ,ll���<цd�I�$cnn�إ����4M��l�����dD��������^�� ��<�N�Z������������(dY~�k�j5���͢�X,��ٹ�~os���V�hp��m��ߏ��[��
�=��hC2"��%�����K��U!""���w"""�9�,�F�������w I<�U>�5���:���D�.���L��,kk�H��z�y�^,..����^S�T����r�S-�9�`ccw�F_�:�e�������%""��$app��cp��)���������0M6��s</m���\�^���
�ł�ɨ4�������#6�9L�����N� """j'vlQOQU����uUݗ^�����dO*������:���D%ܿ�`��Z˲����T��gn�h4������r�^�H$����z��d����0��p�6^�.]�qzz���U$gh4-LIDDD�̲,��T*���4����$IB8���0$IB�T�Dwr��7�H�A�e[Ӂ�S��iJ���	����2*�2b���M�n��`�d�e�)!Q�1M�����a۝�BDDD�.��NDDD�DE1c�楟�����ve��Cǻ���ND=B%,//#
_YkY66�q~�hC2�Ap��8�����4M������ȹ`�Ӣ����55���T�U���SV����P(���;�F#x���t]�������z�}��� ��g�:������[lh��177;�c�l++��)���A�(fMӌ�0�Np'""���(��j�篨����EiW�[�׿�%NOO:���@E,..!�ب�������N�,--app���j��G�"�N9��zU8���"���@U�k_�\.coo�ۛ(l�!""���j5��'�J%!I|>ߕS�?�(��B�,�(�l��+��H���¶�#�B!d27z�V�r	�z�XW5�{<}H�8ɝ��)�eyE�3M�Ng!"""jNp'""���r�&5M۲,K����gf���K$���>�t"jA�hn�F��귶6������X\\���&�Lbss��r�`���B�t�R�����H&�[�����z���������!���5u�F����c�08ѝZK%��΢����z������x�aff�Vm*����
�܉�"���x�T*��NDDD�'�QO�g�i�/��D"����ѵ&j�'5|��h4��BD�Ys{�V�����o���~,..75!��� [[[�,N���	�������DS�-~W>����6vwwP��[�����z����d28;;�i���jt�$	�PCC� �R��&Rj˲�J%�i"����HeY��� �R�)�J�t]G$r�P���ׇT*نdDD=I�,뫦i�/�BDDD�46�ѭ�(�?�u�_\V#^��W��z�����/~���D�c��A���b�K��������c�SQ�����ILNN�n�1kk�����������,&&&�v{�}�l6���u<}��j��DDDԋ�@.����E����F�p8���a ݩ�J�"r�"�($�ꏒA@4���B&����ۨX,�0D"�+k}>�^/R�T���4�UU]5c��Y�������DDDt�)�(fM��]V45=��}����t�%����t:9L����>�|oo����NQ���öה�%����V�:��z����ݻw����U,��<}��b�eو���~�$I;w�:��w��u�������5\.���^S(䱺�M�LF�46v��j�3lll����ZOłi�a |�GDDD�'�ѭ�(ʿ7��j\.^�+�e�]�n�F���>��F����.���5�?y����[������� �^�L�ce�16>Ы��|������|�K�5�^�e��<���5�)����gY��NN�Q��������,ˈD��i�(�K��^c�\.�~{��\.7�P��ٻ�ظ�;O�߳־Wq%R�wI���n/m��n_w?L�y�`���	�� y� @� ��� �� �)q_�=ݶ���u���⾈�ĭX���%�4���U��� �H�w�_@dթs~��?�E�\nqB�l6A����ֺ�n��6$�6$#"�YLӴ)�2h�_t:Q�������z������Ϩ�k�o��Gڔ��=z�+��G;��Zljj��j����a�Q����caa	��X�7M��ϱ����7z?�SS����n����뫈FϸH������4M��7��.��ʍ�P}}}�Vk(-HK7�i�H$��4�@�PspI���ߏJ��|��-zQ:��(����4�{`��lr'"j�4�����iZ��Y����Z��DDD��~nF�H$�|خ<=/=ãG;��Zlrr
CCÖj_�8���~�Q������Դ�&�b�����&b���(
FG�0;;��}��x=�}}}�h��79%Qc�nt/�JW��(
"�>�Ba��%NҦ���e�N�� I�o/��p8EQ�J�ڐ��-�NA�ex������$�g���� �0�_t:Q+������z��(�PӴxY� ��׾��ޮX=�V��o~�#N=%�q��c�m����%�?�kq"�Q133�[�F,��籲��|��ɨ�I��[�F0?� �?`yq�g���bX[[���)4MkzN"""��U(�qrr�J��9��Fw�͆���|~
yT��$���R����>�6���^���d�a�8!�[*�����x�uk}>�@6�!�DD�dƀ��k���w:Q�]�. �u'���6�uY������oW����_�-�vw;��Zhx�&&&-�aww�ŉ�TՆ��K7�_;?�bkk��	�t5� ```��cPU���r��~p��b���|DDDD�$�"����\����    IDAT������s�˥&���FEܽ;���[��)
X]]�n=�������pzz��DDD7�(��0 �Ng!"""j&Np'""���(��������8�N|�+_�(���Ӣ�3<z���1������155+�OOO�����P�vn�����t^����4���{{�0M�_���D�0?����H��.e%	ll�������Q�1M�|��'�V�p�=W:/r�\��fG6��T��4�L&Q.��,��*����fQ��ɽ�$�	�l6x<����P�b�b�Ɉ�n�4튢���~��5܉����8���j�_�N�o}��mJ��4M�'?���&�a�P���nZ���b{{����"���(�&F�j5��=C4mq2�U>������(Wz�T*���5��
u=�4��eqzzM���x� <���!�"��,�ҕ
y$�I�AȲ\�^�$����R��Pȷ!!�S2������S) #�ˡT�nDD�b��o���Q�V������z܉����|b��e�H��Ю<=�ѣ_����1��E�~?-5MD�g���wB�=w�brr�`�y&��������ٴ@�s:]�������v��#�Jacc/_������z�i��f3899�r��(�������l8�+�V�������`��?w�p�("�N�!!�S"����u��o���*�J���<�0��1���t"""�fa�;�UU��V��g�������ׯ�,E�u����_u:�������2$��[�D"���u���������ܺ5b��D"����j�&�^d��099���)S�>_&����:^�8D��F	"""�m����N ����[o�e�P�p�J�R�Q��麎��(�v;�nk��>�^��D�i�8!�S<����ἴNED"}H��\�LD�$�aܶ�l�꺾��,DDDD��w"""��i����yi����F��+SO�u?����Q�r8X^�EQ�֦�)���r[���*�
�,s||���M6(PCDQ­[#��[����XS �E��l���=N $""��0�R)D�g�$	n���FwUU����ߏ|>�Z��{�:�4�ǡi�� ���;N�B!$�Ih�����6�x~���Q����3@D�$�i��i��C�s5܉���'(���u]���j�v;����Z�DL��<}����N� ���lX^���V�6���ٳ�ކd�..�����n+��a����˗/Z��zM$҇��ED"}E���+�
�?����
�Bu]בH$��CUU���o�����@&��a�Y��eQ,�,�߿^X��d�S�X�C0�����J��.��9�-5�i�.UU����;������}5>��������pj�楝�_��0v��ۛ!�J�����8���)��{���|+i (�Jx��wr�1�`sss�$�R}�V���*2�t��Q/�x<�������ŋC�0�c ���z}�{w��\�vn����.����a���D4mq2j'EQq��}8��1
<y��VkC2"��&�b�0��L����/%""��'��_�q���`0�>�����7���O~�#�J�NG!�&�$KK��v���V*<}��
'���۷�`zz�h�rA���ӧOP(�[��z���0>>��������4pvv���gH�R\lGDDDt�J����S��yx<^(����("����j�"w�!k��*��c��}�v��p�  ����^a:��$"�������
�ߏX���ޓi��,����7��BDDD�>��NDDD]�n��^�Z�������|�k��S}��k8<<�t"j2Q���di�_�V�ӧ��Х�����)ܾ}V7{K&x��j5N��A���0�������&b�VW�!�r�(QJ�"NN�Q�T��x�6��:EQ�����#�ϡV�e�O�uD�Q8�\�������B"�`�s��4�T}}}u��l6x<^6�5�i�㊢��a�u:�U��������i�?7M��;$����lW����f��?��#fg�
���꺆���(8��WH�������[>������0M6S}�P��K���(��J�������ch�ւ�DDDD7C>����	4M���m����p`pp6��l���.�4��`� �,tu�\��|H$����Z�L��{.��6�#"�Y� `��?�t"""��b�;u-Y��]���e5���_�]ȲܮX=�4M���� ��w:
5����f�0����l6ۆT���bi��~��z�4����/[��z������<n߾s�s�\.���u�Z�NDDDD�`�&����� I�n���:� ���```���:Y��fP,
� �V���Ba$	�:���J��\.�H���s��邢(H&mJGDԛL�*�rbƣNg!"""�
6�Q�R ��i��eE��?@_�����n��;����t"j���	׭3M�H&�mHE��p8��|.��R}�V���3���'�n�(
&&�055������j��;���A�\nAB""""�u�d�X�Gc�m�$!
!��X,��*H&�������~��).x��r�b�H�n���s��D:�jS:"����4�{ ܚ�����܉���+)��ot]�Y�������M���W,�ӟ~�m��z���wp�Ψ�ڭ�M�b�Dm��z��|6��R}�T�ӧO���Z���]� ���� 4vf�NN�����\�;E�C�V��y�ln���6t������E&����-JJ��Z�";����~T�$�� �ϡT*�!!�Z�XD�VC(�[����i���4UEQa|��Y�����n/"""�:�c�\.��y�~�_���a``�]�z�O>�1���:��������s�j��vqt��ŉ�]"�ff� �����d2���unO�r�ݘ�������D��;(�ٴBD�u11V�,��,ADH�Q� �"$Iz�o�9]��qoE�s_Wu]�i��<M�>���iB�u��և]7`�ƫ3���i��#�V��E�t��ϥ�:pt��s���^�$	33s�Ö�M����&��h��Q�ܾ}ccw-T�X__C,ky&"�^%��r���<�L�������������,ˏ4M�tz���|�+_kW��vxx�O��N� �&��XZZ� �op><<���~RQ;�����^8;;����S�dY��������kN�X�����d�Q�E��@QT(�I�!��$����k�3_^cz73��A�th������4��W���|pw."��,+��9^>����6��L�Q/�{w##�-��Eo���oVV� ��s
�Uɲ�7��}��9�����;W􉈈�F��lT�T��Q���O�b��j���~����NG!�&q�\�w���N$�u''����nC*j���1ܹ3j���TO(���l6[���j5���(�n0A��*Ey��E���__�����$�ӑ{��k�V��iz��_W�|����n&�Ӊ��	��+��aoo�Z��ɨ�p!��6==ciVM����G(�mHEDԛǗK���;������*6�QW�$)��z�e5ss�XZ�׮H=����x�|��1��Il6����R3��y xøۉ����Y��]����~�z&'�>�4M����`��� ]�p1m�fSa�;��*l6TU����p�a��{j�z�2M�Z�J�U�{�R����j�r��w:*�H(���G��j����}��/�]��fg� ��w��T*���U��� A0;;�H��5�r��Ǐr��I�t���X�sYŻDDD�5dY�/5M�g����v|�?��(�ճb�s�����1��IdYƽ{�r���&�	��>�4� �2���-�뺎��U$��'�n$�n߾���ۖOޖJ�����b�ЂtD�n�(��p�nw�n�����i�fS�(j�#R��jUT*U��%��e�J���0�NG$�� ���1::fiG�_��尳��\.ۂt��^/�,_���X]}�f� �"������r9<}������HQ���V�����ADDDd܉���[�DQL�a��苿�%���mW��e����"��t:
5� \�(x��&���X\\���T_�V���S���'�nG011���S��U*����T�'����f��n���x����sUe;5�R�|n���i�D�TU�ݻ���h��׻����C׹��&�Á��e˻��e<{��b��ɨ�$Iƽ{��v���r0�Չ�X0��7 �����c�;uY����i��e5�@�����M�����V:���dff�R��z�n���K����={�J���d�m�v;&'��>�0�xq��/_pj/�5&"l6\.�N'�N�n7$I�t<�!�@�\B�P@�\F�P@�X@�P�a���:��������Kد�V+���E,vނd��TU���<���Z����g�f9��۩�<������[[�mHED�{E��k��?�t"""�z��EDDDמ��)���i������!"��v��Y�\���ǜ�L�#������u�ZO�<�Գ������I�-է�)���B�8A�>kpp��WjpM$���F�\nA2"�
EQ�t^4���a�����t]���r��b��b��R��b��B�M�u:э'���166f���ے����Q��>K�$���#����0ll�#��8����½{ ���S�qxx��PDD=F��r��y�pѵ�;DDDt�ɲ�KM�>���ΝQ|�w�ܮH=�G?��ѳN� �&���t�:�0������u�P(���y��k�ވ�b��\�tm��˅��x�ކ��T*���s	�.�.�.�n�n��bmW�^�iLӄ�k0���0�]�a�4M`�Y����>�~�a0M��>�QK�7/�2A�$IE���O���	�$�3��d�J�B�B�|�B�b�iv:э��6ܽ{���a��0t���%�3A���$���-՛����M���H����X\\�tmckk���DDW ��4M��N� """�܉���Z���_+��?��F�$�鷾}�-������o����ADM
�0?�A�������������~LO�Z�?�p||���] l"�� �֭���Y^$�i�899���s�C�F����r��v�����e����躎Z��j�M�A�t�M�P�ՠ�:4M{����.>��&Y�!�2$I�,Ko}.C�$(�I���)�UU�(
D���9��a(����������8흨�� &'��t:>6��`kk�b�ɨ����Ĥ����]�la"j���>���׭3M��+H&�mHED�[EyP��w:ѻ��"""��$��u}䲚��%,,,�+RϪT*����A�R�t"zO�����9=�m��;8>>jC*j�����6�4M���������kx�>LMM_i�`:����6
6#���f���y��r����>��D�ZE�RE�VE�VC�VC�ZE��ٯk�*wi����e��󷿶�T���~΀j��|>�\��G�j�ӱ�z� ���]K�I�f�&��^��`���������������x�|�ũ��n߾����u�t]Ǔ'����ې���wȲ��i�l�s�܉����R��j����Éo}�mn������88��t"zO���?���oD���02rw�[�5���H$�-NE�B%����֭��'>W�U<��h���5�,�p�\�z}����x<]�dl�j5�J�r�U#{�U�z�R�J�ɝD�;A�(�mxw8��m��T�l��Y;�Z�"�˽i|�f3��N�Dv����C[(����l6ۂdԭ� ��,_>99����kYw������u�j�?D�\nC*"�ޡ��X�V�m�s}6��u%���6�{Y���%�ݭ?Ņ.���G?�A�c�{R��?��Q;�X�������n&`rrCCÖ�k�VWW�$Bo�!LNN�n�7t�i�899���>t]kQ:��C��&�{��x����4Q.�Q.�P*�����j����7������>��p8.>��l/��R��|>�l6���]��N�"�j�P�Wxm3qzz���]��n���KPU���h�[[�\P��A�����p��b��ǏA��>���*Q�a��%"""��E����n$EQ��Z���_V���������I~�����c6<u9Q��|^��nm&����Sn���A�����,�W*e��<E�Xlq2���`bb}}���尽�ɭ߉ރ�n5��b:����u�L�iJ�"J�������r	�J��bd� ���o��v;��?�N'$�z��f�曆�L&�L&�j���XD]G�$ܹs�]���2����J%[�����n��Ҳ��� �H$����k ]�׼��ZKU�Z�V�Y�s���y焈��n:�(�I�0�ˊ���G����>z���U<[y��D�A���B!N��	DQ���<�����b����'�T،E@?��'�(��f���qpp����lh%j� p:��ih���٫�*
���
���Fv�v�e.�N��N�.��������Q�V�ɤ��d��f����]����x<������n��h�{{���j-HF�FUU,..[�Y�d�X]}�k!]LQT<x� v��n��y�mHED�DQ,����DDDt�\�+�DDDD dY���i]V3<<��~��mJԻ
���ݿ���.7>>�[�F��U�U<~��r���dY���|��Sˀ�i�Ϟ=eAUULMM[Z�������P*�ѕ�I���z�4�{�>H���X  �4P(Q*Q,Q,^�Y�K��$I����y���t:��y]vs�4�l�Ք�4��,��.!FFn�ΝQ���б�j;;[���-JG�����"|>���|>����j�'�Vq8��E�[{xx����6�""�����Z��:������m��
0�+6�m�Z�n�����A��?����>z�O>��w:����ALO�ԭ�uO�<B>�oC*j�F'ԥ��t���n�H���SOm�4ϟ�����EɈ�� p�������|7뵂�i(
��s��r((
l����zw��I�.��x<�j���V3M�|�t
�T�L��{D���p`rr�@��cc�s��ls!/AE���!�X�/�KXYy�Ż]���by���E��8?��!Q��p:�ÅB��Y����^c�;]+�,?�4m�����)|��o�+R�::z����N� ��������A����4M��� �L�)5��n���=8����D"���56S�p�,���q5|l"����*�LL�����n�&J�"
��i�\�\�*'���$��w���������S�Б�d�J%�Lz7M�cy�����LLL@�[�Y�V����D���o:A055���AK��j++OP(Z��Z%
c~~��n.�a�����f�mJFD��dY���i_�t"""����NDDD׆�n��r��ח�Ȋ��>�3���v��I����o�u1�ݎ>�4�ykkgg�mHE��t:��t6��R}4����n�`0���i�?7�U�U��n#��(Q��hh��������E��i�(���r�f���s(
|�'�CD��nx<�W^8�κMq��i��4����ߗ�b����)D"֦p�-=���6t]oA2�&���uk�R������3d����V���Tݺj��G��R)�!Q�S�~�V{��DDDD ܉����$酮�ޅX^��ٹ�vE�YO�<���z�c�I������rխ=8����A�CQKx<^,--Y�fxt�{{�-NEי$�����h�{{���j-HF�=TՆ`0�`0�@ ��D��0ߚ�~1�=��sg�&E	�n�^�n�N��#Y��*��$R�R�_��FI���    IDAT���jx�f�\���&��T��Q�Ý;��ju]���
��tkCQ�ܽ;����u���<�<yą0DDȲ��i�l�slp'""�kBU���Z��ߗ�8�N|�oC��v��I�L���w�CԥA���"B�P��X���kmHE�������d�u���x�|�ũ�:�����BCP	��[H��D7� ��|C�p��m�P�T��f�4��r96���,�p�/��{�^x�>�����i"��!�L �J"���.t�Ȳ��w��`���{{�|��.&{O��mp�б���T*��`�ss�D���%�	��>��GDD�l�?�T*��t""""6�ѵ IRR���e5_��/[��C����5Σ�N� �+������pݺl6��O�p1K���|X\\�$I����vqt��ũ躒$	w�[znx�i�8:z���}>WЍ��*� B���vYn�"Z�4Q*��d�|�˥�}"�NUm��|��|�z}�x�h�m�Z��t:�T*�d2�J�Ҷ�M�i�@ SSӰ�W,����l6ۢd����133A���m������ې��MEܻw��n����ކTDD�M��S]�_mHDDD�dlp'""��SU���V���e5�P�G�lW��u����ŧ��ADW400��険u�r�?D�ZmC*j6�Ϗ��%K��i`ss���mHFב�����,����677�ɤ[���z����G0D0���j���u�\�M3{6���km��D�<���绘������x!�b۾>�C2�D"�tw�DQ���FFF��-M���x�|�9o�P(���K��M���cmHFͦ�6<x����̶�7qzzچTDD�MQ���V��/��ADDD7܉����dQ��a\ڕ�{����뫿�(�[�Z�w?���r���A,..՝>��:?~�B!ߦd�L�`��n�����5$��6$��FE���ŭ[������#<����&�5!I����0��Pۦ�_L\N#�I#�� ���4لJԋA���y5����oy��U�V�H��ǑN���K=-bzz�R���
�67ב����M������h�<�4�Wȹ�e7�x<�w�>D���a�4����4{]FŜa>pU-u܉����E��j��?��fxx_���۔�w=|�+�lou:]������X�!kbuu����F�`��֦�i����d2�6$����tbvvn������2��6�N�Z����EA0B$҇@ Ж�ʺ�#��"�J"�N!�˃��n&A�v���^5�� I�_\cR��8�8wr��$I2���188��q�i�ŋC���7������E�[k�&��6���!5[$���BݺZ��Ǐ�T*�!Q�RU���V��U�s���w"""�$� 	�4�y�W|�O�����\='��������#���,+x��8�nt �������6��f�#���� �oĬ�jXYy�)�7T� ����N��u��vv����N��nw �hj���h�%O�0����f^5�g`���LD����@ ����7�i"�;iv/�-�~D��0==Uml�{:����*�J���u�t:��t��. lr�n��c�sg�n]�X����iZ�Cu)Q��a�pEu܉���cdY���i]Vsw|_��o�+R�������u!A����@ P����[[mHE���avv�P�-z�Z���
�6$��DQLO� 
7t\�Z���wv����zGG,-{͢��i�R)�rYډ�q�(������#��q�շi
�<��8���Q,��z�,˘��D�@C�i����-�b�-JFי�n���=����wv�qrr��T�
��s���[�L&���¡0DD�P�_�j����9����fb�;u���U.�M�|��2I���N����z���>��g��ADW099����u�L++O�lׅ���03��v�\ ���l�S*c�slooC�j-JF�^.��H���[��^�V�J%�H$�J%9ّ�ZBQ�W���B��7�X, ���<����"�>LNNAQ�����F7��v��n�\rww��G-NE�&�"������֭=:z����6�""�N� .�k0��s� �܉���#dY�TӴKG����cy�^�"�$M���_|�o\u�[�F0>>Q��\.�ѣ_�Vck������̬���J���O�T�n�7�(������S�U����x<ֺpDm�����p�n��Ŕ�,�8��r�\˾����_5����-�'^�ݩW�����i�Í�tT,����|>ߢdt]�����{p:]����vqt��ũ��TUŃ�f��xl{{��'mHEDԝdY�+M����9�����a�;���(�j�_^V��*>���CU�v��IO�<���z�cQ��� ��6�躎Ǐr�w�����-/��XYy�����tbvvn����b�vv��腺���H����9��e�RI�R)Ni'�kG�$���݃�����b�;��H�SSS�e���M�ċ�888 `�,]?��bi�\.kM��8<<hm(j:�ۍ{�@��K�L����S�ө6%#"�.� ����V*��Ng!""����DDD�v�,oj�6}Y��`zz�]�zR.�����0��Q��N�| I�/�3M��+H&�mJF��hs�ӧ�Q.�[�����a��O@E��h����m��G[���u�N��Z��~1�=�x<�d2�&N"�*n��P�pn��e�'����<���(*�J˾Q+�lv�����4t\2������j���u�(*����rY[T���<���T�l�p���w�V����.@D��,?�4��N� ""����DDD�Vv������.�q�\��G߆(^>Y�.����V%�2�$���,m�������6��f��䔥�b����'l,�AE���B�pC��rYll��F<uYV�D��? ��ג�aR��8�8׈�'�l6�!�Ba���Eq֙�d����q~��0�U��oa||��ߍZ����M$�&��F�e,--���Z�g�{w�}����֭+
x��!t]oC*"��#���h��i�s���w"""j+I�u]�}Y͗��e�mS��tt�?��'��AD��_@8�[wvv����6$�f���w�-�
��<a#�133UU-c�&^�8���L�la:��E�@����#��_���jH&H$H&lP!��&I�� "�B�0d�򝠮��b�h��x���</fg��p8:���{{���a���055�����u�xkk�mHDD�}^��=��DDDtsp,*����_ӴtY���~ؒF��B�u��'?F�M�D]ettCC�u�2�4�������\L��T��籲�S2oA0::���iH����r����g�F�Z���Y��~ܹ3�����r5���T*�����{���E<C�X`&�<�4Q*��qtt�L&]ס���5�� �ӉH�CCC����j\�I�Z�Z���)TU���|���E8A:��{��0�b1��~�l���>��$!�J�!5K2�����~�����a�f3mJFD�=��l�_꺾��,DDDt3�s�����F�s�0.M��o��OR�w[]}��g+��AD��XXX@��h�r	�=�M�.388���K�ln�YE���,�`C��b���ނ�i-JF�N�������,Ԩb��X���9
�B�����y�>D"D"}��lM�b��h���Q���?>Q���LOOC���躎��-��G[���I�����?`���`���EM�(
�������ibuu�d�MɈ���$I/t]���DDDt3p�;���(�X���YM��KK��ԓ��"~����4��2Q�p8�X\\�(^��L�4<y��J�Mɨ�,7�g�Y��<a�������|n���1��cww���a|���I�d`jj
cc����M�  �R''�������>��4�C�RA*����K��)���y��EA ��[����a��wϠk�X,��<
��Swz�k�("���p �L���0M�X^��n4p�)'}w�0�N���? Q�Y'��b�s^�!"�5�i�TU��u��������8������BŴa��j����p�]�z���S�xq��Dd�$I���\�:�&VW�!�H�%5G� fff`�w&���g+�u�8�	FFncl�.��e�\.���u�J�&#�:�ǃ��!���C��;S�\.#��#;G&�""��#���"�C$��6w���i���qrr�|>���&j���[� �������y����\��Ess���]�~�|/_�hq*j�p8���źu�|�?�a�mHED�=$I:�u���9�����q�;�������i߼�f��-��ε+RO��cx��Q�cQfg�,m}�������6$�f�D�033k��9�I�jn��^�(
��144�@s����c���qJ5];�,�� ��3�sg���I���TʈF����.��v�L&��	Q�T*$�I!�NB�u����,PE�CC�o�CK�"�_ӵ��e�L����(��cTU��� ��
�B�R�]Lr���r��t֭���j��rmHG�P,!�"|>��u����#��)Qw0Mӥ(J�0�_v:�6Np'""�V�DQ���λ� ����'��<�󙦉��w�d�ӝ�����w06v�n]<��ڳ6$�f�D�0;;g��}ee���n �ߏ�ٹ���V*elll �I�0Q�~!7�� j��ϣ8?�"��6�q���>A����ߏp8���8t]��y�������N׃$I����PCǝ��`ww�a�(]� b~~�P�R���&NO9��{X\\D0X��www��Gm�DD�=^���t�n"""���	�DDD�R���O��岚��1LLN�+RO����ݝN� "�� ��g�6@�E�����y	�Ø����ܞ�f����{��;wF1==Y�-�����
J�b�Y��6������G�r�؉���@<���s��l!�LpR;Q���%��q�P(@�$����~�=�}pp�HA@�T���(�4�H$P*-/��x<CH���4��)��L�b1��K��C�0��*�yNr��d�H_��� 2�4��r��]�i�TU�u]���Y����wq�;��]Ōa�
DQğ~��p�����S�Z��J�NG!"�v;<����3]����C����[�A��/Zj����x��1"z��(����4�5�4���/_�ha2"��� ��������Z&�F4E,v��B"�kLUU��������nCG4z���#����=.�U8��-4�3��������0]�(bqq��ibss���6$�fp�ܸ�AݝKj�*>���EŒa ��BDDD-�	�DDD�2���K]�\V311��ѱvE�I�VW��-Q��$	���a����nn�#�I�!5C ��B#��O����</������Z>�R��ٳ6�P�I����A���bd�vӦ���e���`kkGG/���8�����u�l��'��bд�v{C;�|A���>44�P( (0M����i��3Ȳ�����(��D�`�ِL� �g�W���$w��W�z� ��(��(8���jU��eD"�K�$I��@4z��*"�WL�TE����BDDD��܉���U܂ �L�|�OI����������<���w�D�%�����խ;<<���~Q3�|>,..ם� ��Es{�VkC2ꔑ����PCp"���>PG9�Nc`` ��~���i����(��3d�٦<&u��@����AD"K�<��V�8==���	'�R����cjj����ײ�,��W�s��$I���|>�Z�4����x<ކd����uk�n]4z��͍6$""��(V_Mq�v:�Np'""��P�_뺾xY����DH�����_ ��t:Y02r�ҍ�d2����6$�f�z}XZ���^,�����^&Ifg�p�ֈ��v�4���!����`�:D@ ���&&&��z�Ҩ���pxx���M��q6|��r��x<���c��e�l6����b:��n݂��}3U���
����~?TU�t��fC� ��f{��$�8� l�˟�A@$A>�G�TjSBz�t
����:�ۍZ��\.צdDDכi���(a�0>�t"""�=��NDDD��!a��;��E�G���7�ݢ�3��?�t"� `qq�n�k�T£G���.��z��t�Rs{�T'�Q����W9��/��rY>�R�`cc��ը#E����`�ۛ��j��NOOQ*��DD�=<���Yn�N �B''ǈFϠ�zS��
Qq��8��oY>�4M��?�˗/Z��:M�e,-݃��[k�VWW�L&ڐ�ޗ,+����?2MO�>A&�nS2"��M��i�~ �DDDDM�	�DDD�t�,�?�a�]V3������vE�9�i�?��S�����n����:VV�p�m��x�XZZ�ԸS*���)��{Y0��ҽ���S��={�b��}��\.�����,��`M$�)���a{{�T�Ɲ*��n�j��d2���c�JE(��ދ�TUE(���0EA�Xd�;��i�H&�(����v��@N��T�i�!)��a��cCu��_Lr#���:n0�L�w����`0�X윯IDD$EQ���;����z'�Q��A87M�W�m6���?��(���Svww�_�]�cQ�(����v��֮��"��!�/�É���CQ�oW_�����c���a##�16v������/qpp �/�>>�##w
���x�j�h''�|�#"�wr8��������zL�D<���Kd��&$$���tbnn��ݚ��<��VQ.�Z��:IQ,/߷�s�����Yl$y~'�oDfD���d�"��M��=�d����/���/��_,`��~X{�Zx�]� �A�yW���FҮ�!Mw��Q���*����}EF�XU��ifd������*���m0����������(�&$���annް.��c}�1����z _숈���p�;])�������iU��z�h̬HC��lⓟ�-��f����۷��H���+���>��f�ݻ� �6��z����56~)�ł��E\�~����F����-���t9�9A�7gLNN��t~�wԑN�qp�Ϟ=};���DDt�fSA6�ś7G(�ː���.\.��q��~(��j���]������l���i�Y�16C�Tb���z7�=
C2�"�"��������r�I���z[���v���l6kR2"��&J�4�i��:6�ѕq���z����b��Á����mm�K�mkk'�ǽ�AD"�(ffn�e�Y<y�gB"�P靈9��F����56�)�Ӊ��{���m��f����r���dD�,+��Ǳ�����1��M�m6�899��������FDD���R)����d �r�>�����@,C,6 (�˜�K]��:���:�`[�\Eтh4M�P(�MHIfSU�t��&w�łp8�T*�E� �����.���|(�˨T*&%#"�_��/� ��BDDDW��DDDte4M�cM�Zvs�޽�p8bV��S�V�٧�B׵^G!���W�5j�67ס��I��,+VW���r�*J��k��9�B���Wa�O����5�����N]g��199�����X���~�R/_������q���J(��L&���#�j5��Z�%I�����!I��
ϻ�kJ�2�4��P[�Z�  ��� ����RU�T���o�ՊP(�d2����f����`�d�� �j���4���:����&"""2�p8��j�C]�/<�p:���o���5v����>�˗/z��ZE��=��ݺZ�4<~��RѤdtY�(bee>��nEQ����S�����$fff���UU����~J)Q�x<LLL"��5M�MӐL&q|��B��1>~�Pz�J�4������5j5���$	���mS�T������C�n{�H    IDAT�cu����o�|����c6D �׋��{�C,����CӸ���F� ���Q �^g!""����2"""�*�iڍVw��G(6)���f�x�՗��AD�ܙE02����E6�1!}A����V�B������ۇ��b���"�]��v���*66֐���F�����۳�y�\.�5�7aoogg����W������j��D"�����
����r��A��������r�P.W�(�'�Q�i�DQ���k�I�066�J��&�!�l6�N��>ɲ�ׇd2]�MJH�Q�ס(��}���ՊL����h�	V�uNӴ?�u"""|lp'""�f�ۧE��h���r�������%G�/>��R��1���h4���ú��#�6!}���9D�Q�:MӰ���b�ӎ�����ݻ�ښ��N:����:��k�� fg�p��4�N�}�|>���gx�t�l��^QJ""�Ω��\.���7��kp8�$���M���µk�p�ݨժh4W��(�͢R� Nx�w�F��u�|ބ�d&EQ��d��v�n��dҤttY�R��p�F�׋J��,D4�t]��r�~WQ��$""��w"""�
?�4m�U���ښhL������l�:��r����lx�\.agg���͛�0>~ͰN�u��l!�͚���������
��x��w_c�ےS�����������JG:����^�z�""�;���T*����\�$��.N���8� EA���>�:�J�T�@�$�q��@  �˅t:��CFQ���F��׈�N'�vR��I�貲�,����x0B*���!D4�]ח4M��^!""���w"""� o��������x��ǜ�~Y�����-���1���	�ֲNUUll�sj� �qc��Sm�>y�ǉkC(��¢���飯�����r2="�(q��u�ךVTU���)vwwq|���DD4��:�3��)��T��^c���Fclt�+�(
����t��^��r��ɤ��ΐ���(�ˈD���Wn��,!�I���.�|ׅ��� /\E~����\�BD#M���.��_s�;}6�ч�SM�Zv ���@��<C���'x��E�cQ��s��u��{��r&$�1>~337۪=8x����.'"3	���������v�T�Z���:��J	��X,���%���C��K�F��7o����d2�f����h�4��i���@�4��.���ns�kt�D"PU�J����(�u�d����j�~�f�!�!��q1���V+�V��D�0z,x<^ @>����LQ4���u�,C��h��F������i�W����b�;]��n��(�o��z�ǋ�>����/��(�䓿E���u"�@<���ú��78<|��@�A��fgg�N#�˗/�32�K��}L:����'aӕE��װ���Xl�$]�{�J%<����,4M�¤DDD���*r�����h4�t:a�^��R�e����(J�
'�Ӈ+�(��Cŋ'=�c�Z��P�T�2�r�� 
������B�`B2��R�����ݲ���V��\�*"]���r�����h�ɐ���.��DDD�!���i7Z<��#��~���ͭM����:]��raqq���� P,���í��\(���b[���������	��,v�w�ޅ��k��������g�0]	A�Ǳ���h4
��z��ɤ���<~��
""Z���X,����r	v�6��R�K�eD"Q6�ӕ�V�H�Rm��#�"��(A��PC�X,B�����A��5�J%��ee��Ba�r���@ �T*	E�ZD4�M�f5M��^!""���w"""���q]Q��-F��|><x���_R�Z�g�~
]g�Q?�X,XY�Yn�@�l6���ΛY}���ayy���zgggx�d߄Td�ߏ������mիj;;[8>>�r2"�(�066�����:����vqx��Z�JS��J�����rYH���y��#�2��"���J����M��\.WۏI���ÁL&�E�C$���j���5^P
�Q*Q�VMHF���:r����-�#���?���S�>���u�6�	�+H����clp'""���cMӦ[<��c�|��~Y�}�L&��Dt���yú��
y�e�\n���mkZr:���� ޘccq,,,�=-�V�acc�<��C�7�/--a|�$I��w�u��vwwpt��F��s�z��D��l��a��H�`���Ze?]��iH$mO� �ۍ@ �L&UU���̒�f�t:�r�[�	��p8�\.�z������TP�U�D[�ɲY��N�LJFD�w��zKӴ���A���h������:�t:������v�χrz�%
y|��罎AD����)ú7oqt�ƄDtY6������Ο������Ɛ33713s���B!���uNƦ
�����k׮@c��D�;;�8==�N!DDD_��=�J�b���r]���fC4C0D�^�y ]Z.�C�ZE(j�h���Ɛ�e�h4LHHfH�Sp�=��oAD8A:��y~+�˰���x<-�<j���IɈ����� � nOBDDDa�;uL���GӴ�V5~��T"�U���/P,z�����������b����]p�w��X�X]���x�c�T���:��	�ł��E����>&�8�����f�ѰX\\���m-��.�����;;�8;;�c����EQ�J�pvvA8��}�Fw;b�1A�jlt��)����r�C�X�o�Z�V�bc�TʨT����H��������-�,B�0���E��l6�P(l��."��"Y��j��4���:6�QG\.�X����h5���Ã�qz�%%	ll��:}�w�F7��M�h6yӪ_	����x�>��j����5ބv������O����qp���+t9�@�������tc{�����;;;H��lr!""�@��D&�A"qA.��n��166�ǋr���Աz��d2�@ ��y�(��D�PU��a]בL�!˶��V�~ ��ߏ�)]ב��06�(�։��@����S�,�h$����; �R������w"""ꈮ��i��V5�<��0+����ӟs*Q����kkw����x�sss��#�u�z��Q��MHE��r���z���zUU�����ӓ.'�a�v{077�7��W.�(
^�~���d�h�v�)���FǻF�����x�Fw�Ӊx|v��R�Ϩ#�fgg�p�\p:�w�`6��Lڄ��m��!�J"
C����6�.��d¤tԩfSA�ZE$mY'I2dYB:��c"I�$I3���a����`�;���vG����@���n�}�1��_��������u"��XSSӆu���qttdB"������fX�(
���Z�����-`ee�����z����u�r�.'�ad��q��Mܾ}�q��wQUGGo����l6�)DDDWHUUd2���/d�x<_�:����k� I2
��Q�Χx'!�"|>�ŀ�ǩ��F:����4�L�h��e���$I\���*�2dY���mY��xP�TP��MJFD�?t]��� p����DDD�6M����iwZ���� ��_��i����F���(D�-v���+-��B�����R�e��㘙i�	���䭭�J%RQ��bcXXX�(�w�P(`cc���c�$�ƍi��/���^j������-��i6�u����f�8;;}۰��DwA��z�/�-��l>��e�Y4u���{N��` �T�Ɲ]��D6�A43����x��:���I�S�\�`6[�ݻ� �T�iR2"��!J�4�i��:6�Q����.ZMow��������Kz��)^�|��D�-� `yy�po��`cc�&oN��P(����6^�t��� �ɘ���kbb�o�i��$�L`{{����Q����	,,,!\�����;;�H�Rll'""2ѻ���,˥�EQD ��X���\�bYjO�TB.�E(��b|��f�!� �ɠ�TLHHݤ(
��"b����N @�V��K��u�lccc-؋��ǃ��3��]���6 ���!6�Q[$I�=UU�Z�ܻw�`ЬHC��lⓟ�-���Ѝӈ��붷�Q,MHD���x��d<� �={���SRQ7	��;wf199��1�^��ӧO8q�:  ���2��H[�1ߦiNOO����d2	U�$N""�^i6�H��8;;�t���jE(F$��(�T�]JKä^�#�J"B�$�z�UB4C��G�^7!!uS�VC�ZC$1���(
�ո�X?j6��ժ�D�-��v;TUE����D4rDI�B�����A��������������u�� \ر����������^� �o��|���3|n{�搿�}�nw`u�n[M������+RQ7Y,,..#m}C�MS�����c�H8���2��qX,֎��4��G���z�==ۉ���ŻF�d2	Y��r9�bS��$I2"�(�~?���Fw���h6�H$���x�p8�-��(��2�Պ		������0~�e� ���d2|^�S�J6���e��@6��""E+���/ �}!��w"""2$I�着��U�ݻ�
�̊4T��:>����4^�!�'V�++�M��r��ۜ�ܧ$I�ݻwa��k���<ybB*�&Y���r~����fS�����L��Ѱp�\��_���T[g�M�u���bgg�$ۉ�����(H&�H�S��m5���@<>�͆B�M�k?]L�4$g�eٰ9 AD$��(�Un��?{o�:Q
��~���rY�Ñ��A�����	�+�H�u�"˲]Uտ�u"""�olp'"""#�?�u����Ӆ�}����~I��H$�z���evv>_�YMӰ���F�����(�XYY��m���簽�����p`u�\.W[��Z��k(�J]NF��j�03s��s�jn�l6���-������h�4$g(�p:]��l/<�ǯAE
������44MC 4��P�$!�ɚ���)����r��t���Z��H$�88�麎B��x|��}I� �2�锉鈈zO������# <)&""�������Z�$韪��k�jVW�!�i�T*����&Q����úgϞ"�Iw?uL,,,��P�T����f������z��f�b����u��.'�A'��q,--��\jQg�P���^�z	Eit!%��V�����Jn����\DQ���G4C��@�R�RR�B�z�P��sP���˅t:�k�.�N#���e^��d�?�>�h4�i��)�ۃj��r��	D4:t]�dYn���7��BDDD���DDDԊ ��t]��n���������hb�����i6���݁��e��L&���g&��Nݾ}�ؘa]�����c4l8d�pKK˰Z�mէ�)lnnBU�]NF�.`qq�xK��*�
�>}���g�ո����hXT*e�^����v|� I"�(�~?J��хJ�
�<��p[�_].|>���z0]בɤ�D����v��v�R� ޏ
�|>��.`�@�d�&�S���u�����s�sQ�b�;]H�����l��V5K�+�F�fE*�b_|�KN�!�#� `yy��S�����'~����'ښ���*66�P�T����ڵ똛�� ��������{�u6{��'�ܹ�����e���E��ϱ���)|DDDC�T*����f^���v����p8���4�Ǥ_U�Ր�d��ZLa�;
��J�x�b����L&�h4f�sw�� �|>gF4�P6����X˟�(��x<8;;31Qo�n�$)�i�/{������܉���B���;]�/�U�e��?�x�i�|����xӁ��LO� ����l�T*���:1;;o�}������D>�7)u���$n޼��Mg��z�ϟt74�Պ�������rw|��6���+��n�����hD躎B!���SX�V��n��#�$��v#��i(��]�J���h �J"A�.�l�=Y��D�ɤ9z�5�M��9�b1�E�~ �j�l����(�ˈ�Z_s����4��%�h�|���?�u"""�O�F#""��d�Z�;UU�U���"��q�"�\.�G���u"��Ϗ;wf_���ȤT�	�Ӊ��ն&�=y��d2iB*ꖛ7o�5� t]���.���t7���8��V:lJ;ol;>>���2�w�!""A��"�N#�L�nw��tvt�(�C�#�Tʨ�j]JJ���l"�8����n7��Z��D���h4&$�n���V��D"0Z�
���f�h��	Gm�V���l�x<-��~?��,�u��h4��$�PӴǽ�BDDD���DDDt�����V�?���j���ih|���P,r"Q��Z�XYY5��V*��������F�$��ރ�v��#�|����L���a|�Z[���b{{�T���hP��n,..�ڵ�m-���l6���M���BӴ.$$""�A�(
�3
y��Ȳ���,cl,�˅|>UU�����iH&p8m�8d�X��P(��0;�*�2TUE0lY'B�0���;�P6�E8i�� ?NOO��|IDW�j��p8�v���z��x�����x�v{�t:a��a�J����A>�u����"""����8*"""	�$�׊���j���zϬHC%�L�g?���AD_����H$ڲF�T|�՗�T*&��v	������������'���3!u�(���_@8i��Ѩcss�R���hY,LM����Ol�'�x��d�鈈�h����8��gT�f���/_����;�Я�qc��]�4M���62�twCQWݼyׯO֕J%��=b�{r�\��!DQlYwvv���]�R�0s8��x<p��p8���j��j��J��b��R�ؕ6��'�z�O���@�w"""�� �T���ʴX,���R7���/>C�\�u"z+�crrʰ��ӧ�f3&$�N���#�e�Y��n�����b�`ii�P���r����ǨV�]NF�(
cyy�`����w�f���(��x����Z+��899� �z=�{���`0�P(�r��	���\�f��T�֏+A�FQ��x;���,�n7�Ng�:Y��p8��)�M����nT�U�G �Kq:��Fc���B4����f��΅� @�e�\.AD����C�F�*a~����\�7#""���w"""����E�oZ�ܺu�S�͠��NN������D��������ԤT*���LJE������Ĥa]�R���zW��P�I���ջ��|m���9ll�CQ�.'�A�p80?�����Z������ۛ�f3��JDDDm�4�l�dv�ð9��dYF<���@>���z�X,�R)#
.��p���X,����Z:�F0��fkY�r� r��Iɨ]�B^���e] @"q�I�D�A199���8\.ץ������v���BaX,��>?�u=(Iҿ�4��E%""�!�w"""�A�BӴG�����گC�e3c�_|�	'����K���z[[l �C�`��s�7��&����hp�� ���X]����V}:����&o �7�������_踡8��������c>������EA"q�B!�����5�ۍx|���A�ޫT*(
�D"���P��l֔|t�t]G:�F45\����9�Oe�Y�bc-�OEQ�����٩�Ɉh��LO� 
����(�p�݈D��e�j��x_Ӵ߽DDD4���NDDD�I�t��l���jnL�`zzƬHC�������:�511�x|ܠJ���o�!�˅���b뷵��c{{����t���{�S��I$ΰ�������pKK+���Z~[�V���>^�8@���RB"""5�Z''�h6��z�m4%�Q�P*y�B �S�l�p��i�>��$!�a�� RU�|�X����#
!�ˡ^��~�i**�
b�X�:���]�1 �    IDAT��B.�33��D.�S��N��p���Z�\��h�6f���OUUy�BDDD ��NDDD_#��h�v�������?���٧?G�V�u"�y���¢a����!NN�MJE�ew�ރ$O;|��)�Ʉ	��y<���k{������������l6��/`jj��|���ի�����"'"""�B����SȲ����ޱ����a�X���ȓ�hԑN������z�p8�N�LHGW��h�Z�"�������d��4)��Z�B�ex<ޖu~��d�&~DtNE\�v��Nl7""�^/|>*��e��A5M��n�#""���w""" 8�IEQ�1��='&'q��S����x�d��1��7���W`��[��E���Ͳ�EE,/���2n�8:z�W�^v?]9�ߏ��UX��ݠ9<|���g]NE�$���2�nO���rYlmm"�J�Q�����NUU�R)�r9x<޶x��o}>b�*�2+EA*�D(n����v��v#�J��w U*e� ��߲�b� ��������ڑ˝���_E��n����������n�͛����z�B�$!A�4T*���u��	�rc����h���������7���jU�����ì<CC�u|��'��H�'��n kY�i��6��{���G(2��f3���5!]�P(���X,�\�����3�~���h08,..���	�bg���:�>}���gP�K	�����[�^���1E���(�mk�J����p8���il`e�f�d�@��N�>��<T.������jY�n��r�_t]G��G<o�Ӥ�n��6Q(LLGD���`f�V[;��� �z���l(�*IҤ�iحlDDD48��NDDD ��u�_����Xl�&F�_�³�O{��p>�l~~��# x���[t�����~��a]�R���:�:P(���R[�<���ɓ}������� �v�:��t:;:V�ua{{�b�K	�����S,pzz
Y��v�\�un�����*�e��"�L����` v�>��d��P&�F0��fkY�p8!�"�٬Iɨ�6����u~��t���FT4��ĤὍ~�p8�v{����>��u}�?��j8"""�{lp'"""H������ڪ棏?���1+���u�~�	��z���<A���Yn}��P����'&��vE"ܾ=kX�(
66�8} E"����5M���	n�M�\KK+���M:�|>���M���rZ%�UU�J������z!IR��Z,D"Qx<^��9���Ť��4MC"�����a��n�#"�Lr����u�L�h��e���C�VC�\2)��P�.Rx7�����dD���q��㽎qi�,��=?7m�C�$ɧi�_t;�76����u]�������&F�^�����^� " ��ӈD�-k4M���:'!��˅����U]ױ���R��M$���b[�TU���&2��	ɨ��������[0�T�m�FO�>���3>�Qߪ�j899������M�t:��C�4�R3�t]G2���nokG �͆`0�T�M�FUU�r9�b1��'�P�\�CY�L>�G<>��^�m�u�|��dD�K��8b��^��`�$�_���9ƪ��� 'R�06��8I��WUU�Uͽ����͊44t]ǧ�~�o�������a3��gϐ�fLJE�Z�X]�Y�k�>}�T*iB*�J�h��m5�(J��k(
&$�~������p8�Q����8>>����E>����h0
y$�	8N8���E�`~��B�f��)���R)X�Vx�>�ZY�!��} 5T���  !�Hp��>�(
t]G lY����ɤ�{!������WF�$�\.�rYÝu]�Z�ֺ�i?7)���� �PE��i�뢯�\.��7�Q��{~p��?�E�c�<Qq��C�\>� r�,���LJE�����`0dX���!w�@�xw�̢���Zk�V��F}�b����[���[.������v"�� �X,E�h��"B����m���zB*�gC���PU��AU5h�MS���fB"�X,�͛�!IRG�i��/��͛7� ��u��4��n�U[.�����&�45u7nL�
y���A�y��?ܽ{>_�C�J_}�%����������Pޟ�f�x��a�(�Mӌo���3!"""j�$I�PQ��iUs��÷�g�	M���?����^G!y7o����-kT��/���zͤTԎ��LNN�e2lmmN}��2>~�o�i��Z�b}}���#���avv�����y�7�x��7��� ��$	�,�j��j��b�~�s��Ͽ�!�V+�w�UU�������|���_�\�ƿ+����OD��j�bf�&���-�������611����m�V*��?f�� ��_@43�;:z�gϞ����e�;���G߹���^�~�/������$I2���`����ԫttt�d�x7VY���F���&D"""�>�w""�f�XNTU���,��?�����?�����D#���au��ᔓ��=�����������lXW�����J���������z�SQ�E7nLcbb�^�*����C�R�N8"�Qa�� �6�l6H����]�$���;߳~7UU�h4�(��M��W�(4����5����Dt	�`�o��n�wt���x��%�i��d�Z��Q�q�� E�����zky]��\�v�n�nY��:���P�.eD�Dܺu�pG�A��:�<�G������by��j{+󈈈h�����hD����_����U���
�����4M�O��(�J��B4�,<��p�o:���ֆI��N���=0lVk6�x��KN0�O\C����Q���077����q����+6m�+�������w�����M�R�c�UUQ��Q���h�����Z���:&}Q��ƍ�~}�pq��e����q1鈊��q���s����}��Y�q��C�l��u��am��ŢIɨ�˫�-k*�
�����C4Db��K��3�j�*���wf�$����p��b�;ш�Z���fs᢯[,V��'����o�Uϟ��_���1�Fޝ;�����&���s���#���?��i4�F���&2��)��jt����F�˩����~�F�L&�'O��^�I�^�Z�p8������?w8��[/@���i�:��j�*��*j���+�
������Ý;�O�T�&prrܥd����☝�E;�����&w.2,^���w!�b˺z����������f�Ç�x���LJED�$�2�����������5V����f��&E"""�>�w""�d�������V5w������fE�����g(�-(Q/���5����F"�0!�kaa	�Hİ����6!]�N��K�66�xc}D��n�����vwt��4ppp����.%#�o��lp:�p8�p:�?�5�w�8���z��j��j��J��>����D>"�� ���	ܸ1�qc��"�}. A�hssm�v7ll��\.�������5ܾ}ǰ.��bcc���}�|ʜA����5�r9S2Q�LO߄���uSi�����ׁA���J���DDD#�w���F��j��f���^�uA�����x��~�٧��A4ҬV+>��p�d2���-�RQ;nܘ���úT*������+3==��ɩ�j��66��l6����� �������TǍ�gg�88x�ED] "����X,��I��nz�wN}'��Ӆ��Yx��5H)���O� ��B�Q�i����cT*��U�����Xܰ���5�??0!�kii�P�eM�V×_~�s+��t�p��l�c�D*�7���X��?n6��eR$"""�lp'""=~AҺ�_8�irr
?��_73�P�u���b��ۉz�Ν9��o�)��/����0)	�BXZZ����J��G������yP��p 
�<666��A.�ss�Om���x�d�L�KɈF��j���������������\�F�b�J�r�R�r '�}���L&���.1�PKm=^���56�Qq��=x<^�Z�x�_dY�ÇC���uGGo���S�R�U�u�6�nO�c�����A�q�NB� 4u]� �������z��DDD#F���S�jU�~�?C(6+��x��%>��^� i~�����vv��L&MHD�p8��!���S`UUţG_�� ������Ͷj��<67�9ml]�v337�xEd"A�r��r��6���v�!Ir������PU��A�T��MӠ�*t][�}����1�7�M��|^���{A ,+A��j� ��X,;*T��R��r��R��r��s�#]������<<������w��d����Q0��b{M��z��Q�VMHFW�f�������|�����G(��&%##�h��U:��#�ϛ����������\�c�T*�ě7�-k$I�g����&E"""�>�w""��"��X�4�vQA$�����af����:��/��|��Q�F�(�x��#8�Ζugg����5)�X,�w�\.�A����M�Ӝ�<(:in�����d�ڈ�e��s[o��m����'O�Jq�Q;A������������jMӠ(
��M�f���~��w��BU��u�f�b�X�6�[a�Xa�Za�Z����}���V�Y�!I,K������T*((�(�(�J�u��`"z?�}zz���������m��A,..���^���c�j�:(|>VW�>�j5<z�%����ED"і5�J_}�ů,�$��699����a�i���Z��)�bE�4�	DDD4D��NDD4BdY����Ъ�����ׯO�ih�~�
�~��^� i337111ٲ�Ѩ�/>��&�Q���9 x��^�z��@t%�]��[�n�U��d���ɛ�#&bvv��ٴ�t:�'O��h4���h�9x<x<^x<�ݞ�lt�4�z�F�Z��x�Į(�ۏ�H]@EH�����݇,�o?l���?�1��J��7��+�����D��\.���v�;:�X,boo��i��Ϗ�啶^��>x�_��͛���677���'$I�Ç��~��%^�|aR*"�P�h��R{ˆ���1��N[�H��E��&E"""�c�;�E1�i������n��G?� ��S�?E.���D��v{p������d2� �/&'�0==cX�N�����7TA<ǝ;�m��ɤ������"�"ffn�ڵ��l6���NN����h0�����������U�u,C���V��V��Ѩ�^����ѨsZ��,��fwY�a��!�2l6�v;�v�@4����b��|>�B��B!�ŭD�"��n`rr��k��������b:�'>��˫m=�W�U��=F�Q7!]���y���ֽ~�
/^<7!�#�`qq�e��k��/Q.�MJED"arr��1���(���j���b����71��׈��F�,��E����V5~�۷�ih��'?��^� Y� �޽�x<-��3����,/�6TT*<z�U˭I�t�ܞN�7��:��G������\��&�f2<y��z��2DV��>��mC��o��5�MT�U�jU�j���W�5��5N@V��v�v�����6��o��jU��y��y
y6{���z1;;����q�TO��s!҈�ɽR�`}�1w[�h��{����akk�tʄTԎ��%�Ñ�5�Bkk�x�M4 ffn����:F�x��%��L�����z��L�DDDD=ԟW������Y,�g��޼��,��?�-X�V3c����l6��D#kbb33>�8�����CQx��Ȳ�>2�RYUU<~���D,6���9�s�!��`kk���GH<>�[�nA۟���Mpj;�6���������&�nS�&*����j�ݟU>ǏA`���t:�t��p8�~�$�׮�F�}�{.��&�4Qq��4&&&��-�F����]d2���h8��}x��vܿ����l⫯�@�V3)�"�2>��{��r�={�]7��� X^^�ۅ�P�V���ײ�j��7�ͻ&E"""�b�;��ey��hl��YXX��*�t����7�_�c�,�Á�?6� ����D�̤TԚ���U�ʝ�-$�I2ч�D���_hkrk>����:TU5!��,˘��C0��\.���=6P�ȑe~ ~ ��v��ב �7���_id��
�I��7��7���r�`��{�y�n>�C6�E.�E�Z�u$"�������f�up��ׯ_����<� ��V�j�+�J��X����{�b�?�.l}���TUŗ_~���D}��v��-��mϞ=A�TjU�����Z��ҤHDDD�#lp'""V���m6���E_E?�͟��4�A����|I�3++w�3�4677LJDF��g099eX���K�|�D�����jn/���`s��C���3ܭ��t]�˗/���k l���g�X��z����xz�G�uT������b�b�SX�+,�����N�n���߿���f�F#�j�p��,"�HG�����pq��XZZn��}}}�&��A;�#���<{�ԄD�^%|�����^��;�|/^<oYc�Z���l�ĤHDDD�#lp'""~nA�_x�azz�����4gg���Y�c��x|w�̶�ᤢ���T�l6���N �pKm6������� ��n`jj
�\z��j���A���^8�>��?{w#I����3s73��-��"2c_2�j����Dt��n�:�B:IЉ��G�B�3$�A I���^+3֌�=c�}���QYU]�0��7w��~W������G�D��y1�K��~�F�F�F�f�V��4vn�^�>�^�~���S��W��F�\B�TB�R�g���=Z����gt}���#��&�I�D��>\���w�g�����S���#OX�q���p�\�⋟X�^s�%���Ph�1&�����8I�B ��#""����:EDDDSIQ��A����j~����v��tc��W�D�i�"��FDUա���~�
�rɦTdF�4lm=�����t������ד.�`mm�J+��v�i����-$�)\�i7��`oo�'�ͣ�*b�8�ݻ���e���!}�����v]�Q��Q,p~~��o����W�f�(��h6���9a�&�`0@��B�RA>����	��NQ����t��:�N畚o?��(��H$��s�.��E��Ѝ�l6��e�i��~F�e��	h��R�n⹹��6Z����AgM�
����x�n
�J%�bq�M*�p�B�.��`0��pĴ.
!���0xM�h������t�;Ƅ�P���
dUU]�9������w""�N��a��O�R��?���t#�E�?���5�D����b1��ZO���7Q'�$I��~�`�|�O�~���S 
css�
�����[ 
cuu훦���xq�irt�Ȳ�{Sڽ^����ah4��k����kh��`�!�4��B �����@ �����n��R��R��r��)�t�|�V�z����}\����VW׆��U�����Ã�S�����>�,���6���w��s:$I'�������rYؔ������d�����0���~ǒe�bF��XDDDd3Np'""��E�[����f5�����]�n�����V��hD��8��{`Z#����NT��H$��u�^�D��5ד���ass{��f�����ln��$I�������c��S�Z;;�P�VF����� �H�޽XZZ���,����||�~��J��L&�w�����H��Q*��l68��n,]�0齌l6����(�h�Zp:��OCt:����H$�s�.B��N'��?�ЍP�TP�V���{�433�o'}���j5�j��YOrw����|���}���}�z=�b1�:UU�(
J��M��L�^��̬�ߢ��C��@��ň �    IDAT�e�I�t*H&����V�$A�h6���!\����u}��hDDDd#6��`�$��B�KGw��~|���pE�j_��q� ���N'66�,o��{��7N'D$ţGK�u�b�^��!}
�ۍ��'�+���jag�)+o8EQ����Tj�N�B���w8::�`���^.��d
,�ѣ%�bqx<���[|�^��R��t�o߾��W���eQ�U��v���n�^��z��B!�����iT�t�] ����"I\.7"�(��� �H��r�0�o��i��t�ɤ�r���J"�2��EA�\���L�V�n�fh��V���ˍB�`O8�h�Fn�š3~ �N۴������p8M�� ��4�/MM�,���v.�k��8�B�?�#�o��K���hl�N�����Y���2��?���./����Ch�fZ�j�pr�ަDdF�4���Zֵ�m<~hC"���ak��Pӈ��6�={�-
7\(�����&Tw:<~�j�:�dD�"!�#�!������S}�P]��Q�V��Jt�^�b��EC��P(�P(��?��"��w��E�{��P(�R�@c$�'Ѩ�T*�ѣ���9���<� ���tF���!�� ����bY�L&1������Or||��g�����2��:�5L��o� ����\Z�i.<x���A�	1���7���C�Tʗ���PQ���~���ш���&��NDDtCɲ��qi��SQ��8�)��h4�_�j�1�n�P(��YT	�������$	[�7� �0����9�p��`{�	�n�em�����SN*��$ܻw��+�5�/��aww�v{�و��$I�ø{����1?�`�2�����t�(
899�˗�89y�R��V�]�G���B��m��e��i����V����A�W:�uN�~ �d
�����.��u:����l6P,
�^�i����&?�P�F�� �HԲ6  ��ʨc�'B�R� ��1m��e�P�L��gc&�@���f���?*�2��M Ms��y�)��R�hZ#��a��M�����F�h#""��|>_������}�h	���6���>�ʥҸc�:�����6E1�;==E&��)�Y\|�D"aY���o'j�dr8���zl9��h�z��kt�<�pS�����M���=��0�|�o޼��Z�
�$!
�Ν�X^^����~����|vv�W�^�ݻ�(h6�lh'1�0�n�P.��N�����z�~�����ǐe^��x��w��^|�b�;M�~��l6Mӆ�� \lOH&��e���7T�^�a�#���P�~�z݆d���>:�6�q�k;��BUU^ۙ �N������TIH�� ���h�TUe��TUE�VE�߿�Fq�� ��""���DDD7��躾q��$��/����k�Z-��_�3�ܿ� �X̴�����`�� ����%˺|>�ׯ_ِ�>�,����B0�������y�N�So�@ ����;|�n�����f����7M�+�����IS��Z��gx��5^�~�B����S"�0�j�P*q~~�t��fBh�f:��c|hvO$�s�.� $IB�����hB
t�]D"��>�!A�JE>�4�Z����!��h4�n��F�aC2�X�f��h��~?:��M>��V�V�L�L��)�
�0P�VmLFD?�t*�F��y�I��^�$EQ"�a��ve""""{������� ����+��ssXZZ�1�Ͱ���B!?�D������ʚ����}�Z-�R�e4ͅ��mˆ����]Ns�`�$auuѨ�$!]`g��ͦ�hfff����s�I��B{{;�t8џ&��`0�;w�|��>�@`4M�N�\�߿�����s�jU�z�k�����躎f��|>���ST*��=8���z���$I�x<��☛������Q6��dj4(���C�M��n$IT�U�z�y�T*8�Nև����:�m��d�r	�h��o<��P(�Nإ����&�H���A�rY�%#�ÁX,>�SA�\(V$W�׮LDDDd6��0N��?�u�?0��⋟\i�&�^_���.E4����x<�5�l'''6%��H����-���ϗa��}�n�M��lyyɤ�Q������A�V�!�M�e<z����=�S�7o^�����D���`~�VVV0?g$M�a�R)����^��۷oP*�j�8��hj]4���e���#�I;������,���!�Hbnn.��� �.��i���}d��\.x��]ot:�H&S��z��}��%�\n��ϒ$!��Z����B�R� ��1}��e�P�L��wǬ�n������^Z#I\.7����Ɉ���H&S�1$I����e���(��xjc4"""16��0�$�+!ĥ;C� �<���H7���Ȥ��At���	ܽ{ϴ���aoo�M�`aa�x²�ŋc�JE��Z\|���9�:!P*�lHEv�4��ۈņ_���v���˛�4q�N�d
>���"����K�^}��`�b������LiO�V�q�%���:���NNNP.���:4M���Yv��`ff333PU�N�Wi�!P(���t�D I�>.��c�4��'n�R���o9�@�$��q�Jen��`�A�v�򚏪�P'��L�j����Y�C	��[��H�D"1��&\.��mI�6��ȦHDDDd6�� ���d0�m��ͭmD"Q�"����?�9o���p`cc˲9�ŋcN�� �P�-[Nx��rx��M��cܻw��`���G��#ND����ز!����vvv�n�F��hx�,#����X^^A,�������� ���ݻ�8>>F>�C����;�[���T*�����F_Yv\����D0���<��dYF���kM�f��R��p8EQ���ߏP(�R�]�G���T(�
�,_eYF<G�X���	�j5��*���i��@��B�մ)�]ס�:�Q�{A�`�t�S���$�3�m�p8��t��\��EQU�_�^�1�܉��nY���aw.{\UU��˟]�������Wx��ݸc�:��D"�5�j�^��)]��tbkkN����v�����4�`��sX\|8T�˗/�N��8����,��և�>+�����p||�`S�_0��������Tj^��� �U4u����ի�x��5���7;��FD��>j�*2�4���7��24�um�G��!�bnn~��a���V�^��L&����;�ϸ\.$I�jUt��'$�\L�/ �BUU�Z�Áh4�B!σ�R)#�B�4Ӻp8�\.��r���"�����t:!�@�R�1}��z�v?\�S�rK�$I���3�"ш��������!�{ ��)}�����9#M?!������D6�z�X^^5m�B`oo�>�>�mee�@д�0��>c�����XYY��G�o�{�''�G�l%�2��Wp������z�.vww��fF��Ȝ��D2����*�޽���{[�&���q|��߿G�Z�w"�`0@�^C6����Z�&$I���fwI���x�H$133UU��t����ꢱ��Q9���ὼ���hؐ��`��b���Z���mc47SL��F�2�ɔ�gmY������r�۸5��R3����` �|���@UU����UUQ�V1\�z%�����"""���DDD7��(����=.I~���f9-�~���	^�|1�D�����n�i���	r9�(���Yܽ{ϲ����RɆD�1�� 677!I�͠��gx�����N��akk������V���y�V�5�dDf$��a,,,byy�X�Z��|��~�w�ޢR��a��>�ah6��#ivw8����G4 �Z-nP����j�T*�D�p8�oIJ��h4�ۍR����B�u
y��q�-Q��""�����P�� �N�x´��r�0t�jU��я��zPU~�Қ��xp��~B�b�qǘ*�,�Z5}o�UUUu]���DDDD��w""���_!.�昛��Ç���s#��_��f���R���ϛ�t�]��f�y<lllX6E
y�y�ڦTtUn���O,  �����ȆTd�P(���'WZ�|~~����:�}�~��avv��k�����뽖�P໦�/����I�Dt����~~~�f�z��5MC4����n7��.7O�Xt���y�!h�6���|>��a�JE�>�d]�Q,��H$,;�\.x<�����U�Z-�\.�|~ӺP(�R��^���ƩZ�"��1��s��h�Zh��6&#��`�h46�A@��r�Q,M��!ք��XDDD4"��DDDt(������|������e��;ѭ�t*��ش��{t��&W���,���܆��L��.vww�^|B)����'C5���% ����$�����:��E3���޿�.��$IB,���C,--!�u0g�vgg�x���ۦ�~�M�Dd��7�����v�Pe�f`3�,���cvv�H��Zm&[�� �l��}}R�\H$��T*<�qC}T*U$IȲ�Ay���CF�\�)]U�RF,��(��H��P(�L&���1�@�߷���ɤy��fn��r�-}G�$�nzH�VU�����BDD4���NDDtH��WB��e���~<y���M5�-~�_��`-��>|�`0dZS.�8|,,,�>U`�ӟ&�,;�����gY[�U���˛�7�$IXXX����П��.��vP,G���;��bnn++k����f������sx��%^�z�j�M�D4t]G�^C:�F>��`0��i����0�}~~.��v��}d!��z�"��P�A�N'��$Z�&Z-nX�	z�.j�����@0�`0@�^�)]��z�T���T���{�5��B!�\�7�:Ȳ�r�dc2"B ��/��˅B!oZ#IҺa�ئHDDD4"lp'""�r��=�����Y����M��}�JO��ݸc�*~�KKK0kZ3{{�؄1N�p�-Yֽ��LچDtU�$a}}�pز��lbg�)t]�!���p`mm����?S�V���Ed�ߏ��`ee�H�Z����R���o�����B�N���F��G�R���)J�"À���xe��T���Y�!��v���d�F��J��H$:��,�H$��$	�Jņ�4j�N�v�xV���_�&T�׃aX7f��~�Z-@�F����Y�	~���HDd�^��X,n�݄��p8�n���^~M�0�����_�A��hDDDt���NDD4�$I�3�0]�����O���O��y�<��w�iFd+	�4�iջwo-'s�h)����ǖ�+�zϟؔ���ѣ%$�I˺^��gϞ���͛B�4lm=F(d�-����s����,ˈ��X^^������ײ��^����=���#�I�X#>=0��z�J���NQ��!I<�'�NJp�݈�H&��e�v�[{h��.r�����u�B�<J�"�����k�Z����F��u�$!��R����ڔ���V�!��|28pqX!��A�6%����p8���H���ǁD6s8Cm٤�8����$I�a�+�2��c��ts!�g���?XX�ݻ�l�4���~��_�f�����133kZ�n�����6�lmm~�ߴF�u��<C��I���޽��s�e������n�@ ���ǖ������x��݈��m�r�q��=���!�L��f������ϟ?���{��56lэ �@��B>���y�^.���|ҿ�t*�#������F����V)]ב�f�t:���ׇp8�b�����iW�׿y�/o�>4��P(��oBU*e$�)�a��d�Y��U�5$�I�Y.��n�F��dD�[��A<���C����i(�KV9
!��]�����������h����_����j~���D���������PU���+8���j��v����1?ǲ����JنDtU�D�-Y�	!����Z�\o�d2���ӛ����t������$$�O���������e�!��^�(�+x��5���P.�1pB$�\���V�����R ��x,�[��$	>���s�#�u�i�J�z�"��PM]��B<G�R���\.���XN�u8�F���r<�0�.�+�H$�u.��a�Z嵆qB���"7��� 2�4	��0���\�~�����k�>&�p*��7��6F"""�k�w""����B�K����q��oؙg�|���[��'�k��Ѳ崶|>���9Ax�</��7,��<޾}mS*��P(������F����P�ې��p��<|�h�)P�Z�����'��IB4���
<X�����	e�n��9�??���)Z��5e%"��^�bggg�t:p:�On�q�\��H$� �f�ɍZ4�F�J�h�t�N��d2�f��7@�XD ���t*�B��r|-�@�V��Yn��B(�K�v�6%�j�Z���x<��88�N�E��n�~�ht�1����B��7�\ IҚ⿳1]#6�M)EQ�۬������t#�|q����q� �5B���躎��<#Y����M�L��.vww8�iy�^lmm�,���k���ِ�F��p`mm���C�L.�����^ӵs8������fg�>���0��y�z�/_�D�\��- !4ud2i� ���iS�EA$���,��'(ӵ�v�(���Pղ^�e��	���SSO�X, �AU͟{M�����}sB����q(�ri�$I���d�<�0F�z33�����~�7[6x���~�@`��AtA�et�]�!B������z��hDDDtM��NDD4�dY��0�]������䧟<�6B�_��^o�Q�nI����iy����7(�J6������X,nZ#������M MӰ����o ��s�~�ʆT4j��ak�1BCvx��^�z�&�V���Ν�X[[C,��yy��0z�.NOOqx��l6�N�sMI��n�^��R����S��m�\�>^��p 
a~~n��v�~��m7��e���-�y���TUE�����0�JE$I˃��N��׊&��Z33)����@Q�ob���dY��f ���#�Nۖ��3�Px�1��0�'�$=0��m�DDDD׈�DDD��%��� .�����T*ec��wzz�W/_�;ѭ1;;�Tjƴ��j���C�я	�XZZ`~`���w�f3����9lm=6];�A�X�����z��=��\l�8<<@:}>�dt�x<^,.>���
B�0d��.C��%�~�/^�R)s[�!�l6�N��R���p���|�PI����0;;�?�n��n��]�z��\.Y����? �ׇb��ÚSl0�R)#�LYn��u�Zͦt4�^���#�u~��F�t�.�V�VC"�0���i:�6�͆�Ɉn�n��H$:�N��(
j����[!��?��IDDDS��������������w��$�˟���I�w��W�D����Dvp:�X_ߴ�P{pp�N�7����p`ss����^��1z"IX[[j�w�^���Fo�P(������z]��>C�Rq2�-|>���|>�'m�������qzz���DDנ�� ��#�>G���v���x<H�fG����щ�M�\F��C$����A$F�P�a�6$�Q��z��jH&��{$F�������j���B�02��E���Vɤ���@ �t:!�<�A�$���qǘ*�$�Z����N��mƿ�+]6�M!!�_!.�:<?��iꕊE���;ѭ����a�U��l��'6%���ђ��-]ױ���tB
����"ff̷$ @�����SR�(��q��o=��h�ٳ�l�k���2���}Rc{��»wo���!
�<�c��F�b�qggg���Pղь��B"�D,�ah��ט�n�F��Z��h4f9���4��Q*�0��ô�t:h�;��������?/N�r��T*e����p���P(�mLF�����s��    IDAT����z/����`<�=:�b��P�}肦�P(L�H��*���6�"""�k�w""�)�r��z���O�j�|��~�]�n����LO��5q��XYY5m|�u{{��uN]�p8��Y�?G�R�!]E2����a�~������t:6��Q������
$i��_�|{{�l��O�D���������|¿$P,���^�~�z�!ĵ�$"�˵�-d�
8x���>���*b�8��8t}��t��:�
�<���P�*�N�D�Z�n׆�4
�f�$Yn$�e�H�\���'���h�[H$��u^��V��cT�U1;;kz=�� ��r8��P���	�>I�0�M�
!���k�0�l�FDDD���DDD��/Ø��A�χ�>���&&�6�f��ͯ����X]]��c~q�ݻ�(�J6%�r:���ڂ��4�+
x��M�hX�`kk��������M�h$I£GK�w�>��>�������1׋�'�������;w���r}��dr�,qvv�7DDc���P(�N�a�^�Лa~HQ.ݓ� ��l��}��`�\.�?0Ԧ�ÁD"�v��mS�R�@UU���:�Ӊ`0�\.�י	�j��r����	���f3t1&��C�e�%�$A�4��Od�n�b�;��OӬ7�Ȳ�h�?�)]6�M���O`ҽ����D"ac�鷷��b�0�D�B8����5�Nϟ��---#4���������	i��ra{���� 8<�G�̃$�L�X__��q̊a8<<���鈓��%!O`}}ss��4���~�����8<<@.�E��mDD�B�uT*���������59��8�ND"Q�R30�F ����}8�i�e�,pь�����Q��mHH�P.�Xl�4\.
��;q*�
�ɤ�u
���ǃ\.gc2��Z��T��y�z��V+<�Ld]���x>i��m�t:�h4���.�B���pє`�;�Q�Ot]����$	_~��}��6���꫟�08��h�$I���&TU5�;:z�f���%�aaaѲ���M��p`{��P7>޾}���sRѨ(����-�Ñ�����vP*G��n�p8�mc������i��x��-�?�J����DDL�z����34u(�:����t:�^4�!8ѝ>Z�X�aC}�$	�h���T*ې�F�P("�Y^O��|B�Z�ڔ��!���T��`���A���5�1B�� ����|~d2i�R�n�~�ht�1��$ɨV+f%�������ƮLDDD�i��NDD4]���Ү�;w�baѺ)�����N1%���ܼ�ͬJ��7o^۔�~�av��W�l6����ٔ��#a}}�r�> ��9�|�L4*.��?jr%p��ٳ�y(�>J4���:�޽U����J/_�����klj$"�2�v�l�r	������d��>LtO&�����jUt�D�1H���a ���E�X�g�)$��R��d2ey�"��j���k�$�t:PU~��.
#��B׹-p������UU��v�h4lLFt;��=A5�����aH�B��ƮLDDD�i��NDD4%4M����o��|����|vE����/��v����s:��oX܈88�7]!I�����@��fc�����.'�N��ŇH�f,���:�����1��� ?~MnEq����g_s�8]Y0����޽M����j�����x�����5&$"�q�v���s�岐e>�o��r:�bq$�)��f��rt5�F�z�X�,[�{�^A
y~�B�� �Z�d��5'��\.���5�IR�T�H$L5eY���E6��1}_����̬iM @:��A"a5Є.H������§(ʿ6���hDDD����NDD4%$I��0�.{�����g��M�����/�����VX\|�P��Bl:�F:}nS"��D"�{�X�p��I�f��`�����bg�)���hB�����t7��\.cww��9]�Ec�*��_0��gN�X,���C���,��n��`�b��l6I�>��݉h4�x<]�9u����n�X, ���tZֻ�n��
y6fN�n��n��X,fZ'I��(��'�O!��:R�������F��C��d���v�v{L)9H��r�lc2�۩�� �A���5,U�P(�MkdY^0������>?M��Oa��ymm�x��H�﷿�Wi����byy��敮�����c�(
67�,W}������ԦT4�`0���u�f"�0����V˦dtݢ�666-�N?�d28<�g����cee,��rԿ!�@6������N95���(�J�dҐ$	^�o�i�?�(ݣ����~����>����0TU���4�h�b�� �P�р��D 4�s8�C�f���?A��.�A��/
#��a0ؔ���^�aff���<�#���@=�d���?�S��t�Ѩ�n
B��_��S""�	�w""�)�(����.{\�e���?jR]��k��w�w�[aee�Ǵ�͛ל�3F��k���5�N��{�1<A\.����z�88�G�R�%]�d2��յ���NN��������B�\X\\�����ml7��eqp��L&�~�MDD����(�KH��a|>�GM�TU�d
�H�v�.K�5]ב����@��@E�Tbs�*����}�ך4M���A>��)�Z�"��H�e>��L��d��$	�P��I��i.�}٠��"Op��H��j��Z��t:ۆa�[�2��a�;�t�s!ĥW��ܽ���3�vw��T*�;э��p��}Ӛv�����l��T*��w�YT	���q��q8x�����7^�~�L&mC*���y,--uK�/�qr�ކd4�E���"VWW�9�t���a�����f���HDD0�J��g�u~���&�k����^/��cȒa��sp���z}��N��x�J�t�'M�b��h4f9�����U��H�Z����Y��.��A�z��t�A�^C2�2���xP��x��h�À��������B�X0�l)IҲ⿵1}6�M8���3]���Y��_��P7n�B���/��D��$I���E1�;::D�ղ)}��i��زl89==E:}nS*���:B��e]6���ׯlHD�p��],.>�0�Ǻ�c���Ȓ,;0?kk�B5L�L{����u}I��h�	!P�Vq~~��` �?�Q��^���s�4�z��9dJ�B!���a��K��D�Z�nǆ�t]�0P*�L&�p�����h6���4Az��P��P�B���@�^��x<aZ���y͐��A�hl�1��$I���h����!�����뼘JDD4���NDD4�dY�s�0.������gvF�z/^���l�1�n�;w� �H�֔�e�}�ƦD�Ckk��Z��9a�ܻwsss�u�Z��ݔ�$	KK�ClW��������ju��h�I����Ylll"�T���\����f3l2$""K&�~J��$I���������D�V�Z@��T*�u�HĲV�e$I4�N!�2�� �Z�D���f4E��g���V��S�%I���C&��1}�j5�M�*��^��z�nc2�ۧ��#Z�飯�B!oZ#I�]�0��M�����#�����h��B����w�V����m�4݄�꫟����D#�(*���M�������1I&��sǪyV`�'�M�p8���e˛��NϞ=��lJF�E�d���!�LU�\?5�HD�Ű���Tj�r��B ����`�L�_[���j>4�g2i ���r��,��H�f��:���(��Q������,�?I��x<�n��F��WӤ����"3�>.�2����,�L�j����ӿQ�˅~����h40;;��r�` �L�s�FL�`�zC]p:������M�?B� �CDD4���NDD4�TU�/u]����$	?��g<�gg�x��Ÿc�x����[��sN`EQ���i�����{>G��rakk��y�u;;���p�഑e�7ӵ�[9�j�����<�B��x<XYYŽ{�?�;�@>����>2�4ۉ����r��t� ���-����p �!O��is�6]��l��h ����Š�:j��M	�:4�8�A�:EQ��x���lJFV>��æu�P��Ƥ����r���_Z#�H��r�dc2�ۧ�� �A���5,I�P�V.}\�P%oƯm�EDDDW�O>DDD��υ�^9������C;�L����7��E4bn���+�7�����8�gL��W���m��8<<�^2	������� pp�oz�&������6B!����5��<E�[i�G(���ŇX^^������P(`��g�m����ׇF�L&����w�FwEQ�L����P��y�~T��B�VC<jk@$ ~��2�r~������jզdd�Z�!�^�e��\��d�A�^����k���G6��{1ш9N�|�qǘ���P(�no�$iY�l�EDDDW�w""�	����`0���j�<��@��HS�V���׿w�oyy^�״���W�Tx�x"�(Mk���}�n�kS*����6T��۷o���I��Cs����*�
vwwx���$aff���BWn�Z��������v�"Ѩ躎b��|>UU-�K��ǋ��9(��j�f��B�S��A�\B,�܈ �P��rنtt]��"b�E5��C�����0A��fffM������m4�M��o&�K���%I��8Q(�Ftu��㉏��sI�����V�ui�"�r���`0�?""�	�w""�	%I��jƣ�w����~W����R�8�D7����,�j�pt�ܦD�}���[p:��u''�9k�ܽ{ss�u�b/^��!]'EQ���c�u��W,�����jv�}�p�뛘���q�Z�^�8ƫW/��vF�����r�~�|�R	n�g��E�O�$����04�%�i���P,��-�@0���D�\�!]!*�2�ɔŴ~	�h�B���'ć�Qf� 
��ɤ�rj�:�$E�����X,r�������=�(SCQ��o$IJ��W6E"""�+`�;���'B�K�,-� �Jٙg��}����o�[]]���ztth:1�Fgq����/�n�qx�!�M��L8���偶v������MUU���^�p������I����`ee��?���O��1�n�_�����!���z]d�4�|>�I�?�p8�D�D�j5���~O��G��G45m�� BUU̘"�~�v�DҴN�e�B!d�Y~���Z�h��]Z�p8��*����@��C<�0���r�84�h��"��cL��-O�Cm�׮LDDD4<6�M EQ������Y�O�%T����^�~��ӓq� �Ѣ��޽gZS�V���k���<z�l�(}x��5���rak��$f]ױ���;S��v�P�gg�8>>q*�&����{������s��ugg�88�G�VAB""���n�p~~�V�	�?0�����4���^/��*t��o��`0@.�G8�p����i(9�}Z�Z-Ȳ�`0dZ��*\.
��M��J�^��̬�+�χz��kWc�j5�D�i�oYq�ݨժ�t��hTz�B��N��ztA�z��k_BUU�g��s�0фa�;��e������d2��;#M�_��+t���J4*�$amm�������p�@�dlnnY>?��9��NmJEfdY���6�n�u�ϟ�R�ؐ�������񓡛�ON��ի�#NE�$�css�h����	!p~~���=�N�$"���j5�N��0Ȳ|���z�����ah4�#JI��0t�rY�����s��~x<n��=-*�
?�n��\^��������zp8��u�`�L��eƠ�n#��1��z}H��6%"��$毕��KC>�3��$�a��M����hHlp'""�<Q!��pi����6B!�	4��\6������FK�f033kZ���IaL�߿o�B��&���.ð)�Y^^j�����x(aʸ\���4� ���89y?�\4�n7VW�p���+O��r����]d�����B�Z�"�I��t���]逗,ˈD��Fch6�<tM .~����~�&h�a��b��4)����P�	��p�Z�'�O�j��D"i��9�NȲ�r�����vL_7UUE��D�ٴ1����t�ů|��e�N�t��"� ������,�����h�(��u]���WU?��Oy��
�>��Zu�1�n,Y����i�h'�����}^������ʚe���h46�"3��wp��]˺R����#�uq�\��~���u�!p|������{�{������{�o�[x��o޼�{1M-]�Q,Q,��z��L�}��bffn��j����&�<�^�P��|><
6�O�0P���L�L��K��H$�\.]ؘ�~��f�rJx @�\桥1h6���5�����N�s�>ш!�����!	�e���(IUU�����+Yc�;���gB�KGz.,>��ܼ�y�Z���o~�+^H%�;w�"��֤���f36%��H��؄�e>):���ݻ��D"S~ kk�:�vw�A�u��ѧ�x<Wjn?:z��Mp1Qrcc�x�J�j`0���78:z�f������f��z�d2h4�W�j���033�0P��G����@������볬�z����(����I�$��'����������f�[FV�W���9��:H��@:��1FLӃ$���#Z��a�@	���yKUWel[Fd���龎��U��f�U��|?T��_��R��n���~�,�7>�n�Fcc�[�� �� >���j��t:���L���~\__�ϙ���.\.����3%IB��E�Z�1����v,���'��"��C�M��/��gve""""klp'""z@$I�cM�������\.�FE�d�n2�Q� z�$I���D��GMӰ���F����D29nZ����������$	���,ק뺎���\����6��������a�͛]���ؐ�2Uubyy��s��~�0\__aww�b��WDD�$5�\__�0t��~���Eсp8�p8�j��n�3Ĥ�����M�n�>���F��݌��p8,���M�����!&EQ`�咍� ��*���M_{}>?���`ܘB4�^>����:ʣ�i=��a�E�?4M�Y""���DDD�(�����3��BX�xic��M�u���z=��%���C�5��g���6%�;N����k����7���5��~˺��=�E�}�x�x�ꋁn6����]�r9���% ������@V?V,����t:]g#=mw���L��4���TՉdr�(�R)�Y�����7��\lrL���~����?�z��F�aS2�G�u��-�b����� r��ݮM��h"I������0P*�#Ѱ��`08������f�{�AH��������,�������p�� �v"���!���q;??���ɨc=YN���+�oM�����'�����<�iM�T�۷G6%"3��SH�&,����pqqaC"�w��in�����|���ϙ�����:��S��~������''�l� "�gG�4�rY�J%�|�Ϛd)� �����h�ZCLJ].���(����6�����H
��� I�ۑ��0��,��< �F^�nw��[� ���!�Nۘ���)���8��-'~��L��#����n!�}�5����p�V���1��4kƟؕ����̱����聐$�?�u���{\����t%'��7_��z}�1�����E�|>Ӛ����T�6%�;ccqLMM��躆��-ް} � ��WM� @�T����M��r�\x�����5���Pඋ�JLNNauu�r������K���Z�)!���n�p}}�n��@ �Y�>�,#�H��r�T*s�3V(�!��@�\.<r���Iś    IDAT��u�r	�D���(��d�<�� ��e$�I��窪��i�V�ژ��^'C�p�A�p8�ݓh���� ������Y�!)��VӴ-#Qlp'""z A�_��{|bb/�����U+|�ݷ��A�dy<^,.. �C��j���  o��ᐰ�����@���)o.= �$���MȲ��N����-h$<���_@QT�ZMӰ���R�hC2z��^/666�',��X�\���և�6�ݩV+H��P��~�^/����Ɛ�CW( I���e������6�G�����"1ߒ��*$IB�P�)��iz���s�N���n�Z��D"a:����"��r�ѐt:mD��Ͼ��\���r�� ���cQlp'""z �n�x����f5/7_tC�n�����-/���r���^�ٔ����͙NN�Z��I�����u�M����]�<=�����PU�e-�۟7Qt`v���V��և!�������GG��vM�*=[��!�ˡ\.���[*�>�ÁXl>��r	�Ɔ��X,@�A�Z���ۍ\��#�Z�
��ey������lrC�P�UM�]��Y�yO�f�a���!����� ���1��i<�@�"��wR��F���[c���m[0"""�Ilp'""z�{]׿������������t]��~��x�hH�� fg_��T��}{lS"���x���l�zavv������MO� ���{����k�/��N�z��N�J�^�ۯMW��������H$���\]]agg�rih������V��t��a��|�k���F"�@��A����Q�T��&wUU�`��ED�QȲbZ���q��CP���L����z}(�Kh�Z6&�z��h4
E����v{P*�n�z$�0�n9�>q8$
��mEQ$M���2�Oc�;������;~dn~��);�<j�߿��w�F���Z]]��4����7�l'`}}ݲ�����LڦL�O0�<�  �R��6��_BUUln~a:Q�N�����kT���C�pHXXX��ܼ�
��R�հ�����+�>��DDDO�a(�K�fo�v�z�vG�Fc���(����}N���냢(VMS4bw��A�['�"����C24:�^ 
�L�|>��9$�n�v�xܴ��rs�ѐt:D"Q8l��{������a��]�������шɲ�74M�O�j~�����o���_��Fc�1���h4���IӚB!����6%�;�d���5�v{{��);b��`ssӲ����`k�5h������n�ZMӰ���J��۟�@ ���Mˆ��uggﱿ��6���^�L�F�`賚��n7��q�z=�j�!����T*AE�M�>��,�P(ؐ�~�n��V��X,fZ�(
EA>�C�V�T��A��5�����R�r;5�MA��XN��j�f��dDχ����u�GC�4�M�a�E��4M�j""�b�;ш����t]���x ��˗vFz�*�2^�ݨc=Y++k��f{{��t:�e"@�d��oX6g�A�^�)���I�V7������G@�eln~��cY��vv�P.�lHF�(���}���%�F��R.�����l6�������K�Q���5dY��7x#�(��D����L�JE8�Z��I�P,���!���p:����}>Z�����pd�F�DҴ* �I�w���:��q��ۃ��+�=/�v�X�rc(ݒe�\ִF�1]��w�"�O`�;���S�0��p]]]E4j>E�>����4�!��ƐJ�O�d2���M
���/Z�`/
x��ԦD���̬�X x���LچD�K|^s����m�JlnN�~?666�F~�������-����v������u�|�j�`�r�����n$I�ZMn|f��"E��緬��p8(�6$���X, �Zt B�0r�ߟ�X�Ղ��1�.�"TU�pP����t��?7���V�r�;����UUG�Q�$	�j��u}�0�`W&"""����NDD4B�,�����;����?�$}ޤ��J�4�����Y��@���A����3��;��z6&#�Ϗ���5N�6�n��`0���eX5�
y��~6I�����^�e������fc�3r7�}qqٲQ����<vv��煈��&�fWW�E~�੗���<J�t]rRz(
��@S���I҆a�\.ې�~��秄D"	Q�։��`0�t����J�T���L��>_��*��V��0>�2}-�w���u�Ph�1�J��{4�0UU��4�뉈�F��DDD#$���u=���T*���;#=j�߽����Q� z����O��\__��&cS"n������Oey�����M��H���/7-���mlo�����C&�"66^�﷞�h:��vQ(p��s��x�����Bw:���-l��0�E�E~���?��x�'�l6�lr��s����r9:�
����P�VlHF?G��E��D,6fZ�(
dY���4�a ����~\__�@��z��� EQP�׹�h:�6"�(��BUU�rY��	A�t]�Kc���]����G0��r���������=��(Jt�>Mo�ߘ���lȳW*5�D"iZ�l6���Ǜy#������5�0��l��w{�d����t��9}��r9�EA���VVV?{t:���������F��n#��� ���5�}l,EQP*��뙸mrw��nr��h6���6$���ѨCUU�|��}>?j���X�ZE$5ݘ%���	�d�z��T�|���������$I���!&�f�V�o�a) 
�뚈��F��DDD#�(��iڿn�8���7�k6�R���ף�A�$%I$��Mԗ��f��i'EQ���n�:�����#�L&155mYwzz�����'`ee�h̲�0��A6���9PUkkH$��=�}��g�u�'#""z�@�TD>���0m��1�ϏXl�J�Ng�)���sp���x<�����*�ͦ-����ED"�My�P�L��F�V�}�f��3�����z��}���^�Uu�Q�F��ݷN�m���>E�bѴD�圮뿷+}�w""����a��:33���I;�<j{�;����	����5H����=�Գ���|>�iM6{����6%���v����ay!�����ȦT�s��/X�n�����&cC*�X,����p����~(�����j�ڐ��/��t�ɤ!�"�~����dYF29AP*�����\.����mZ'b���2����Bit��$	����^��?�R�ӆ���ۿ�Z��n~>�Y�j=����r�;�h�������+EQQ(�MO���B��lc,"""��#a���F��rMi�fڽ>33kW�GO�5��n�1���D"	��eZsyy�N�mS"�@ ����i��ix��ئD�SA���*���v�6���kv�R��*���E��X]]7=�c�^��{���E��bB"""��t]���[|�ݷh6ߌ%��g����$hz�����.
��e�(�X_߀��!��f���u�PP3jo߾��\��FmJD����k��u�ˍ�1N�&� C�5��-ۓ������܉��F@�����~���|��O�z��������c=9� buu�$���4{{{�uNo�� ���x	Y6o�<==A�h}s���ŋ��5����z�+��Tj��/�=>>���K��������#��}�B[[[�T8͕���1i�۸���(�� �f�r��H$�h4>�A��0��e�t:MkEQD,6�|>��T�^����k~!�Pȣ��ؔ�~L�u�z=D"��@ ���0ædT��Mq�?s��������TD�C��F4�(�%l�,!�ϙ��,;u]����DDDD��n���h4��0��w:��H$���}�Wߠ^��:ѓ3>>�x�|J��ŹՅ?�g��������:'��X0���a���s6C?p�x��K�������E#�JM`uu���=�^��Gx����CaDDD��a(�(�������8����r�P,�\���6��G�(�������?|���"b���Ϻ ��H��8=J�Z�p��c�� �R�hW�gO�4Ȳ�?зF�e�Z-�j��Ct�$I�Ƙɲ�R��^�׷F��0���XDDD��qY"""
Y���u=hV3==mW�G�^���&3�DO�(���2�]���p~�FN;ɲb�� ���!o���$IX^^�ln�ժ8=���,�bii�4�_^^�����C�Ȩ����/0?�`:���
�����<�BDD�D��e|���H��?�������W�x<CJFA�����wh4�'������́K��4MÛ7{��W\.���mJE?�����s511i�a�����{�C<��3�������G�Q	�B��k��PUuѦ8DDD�'��Lſ�u���P(���;#=j�opss3�DON*5�Xl̴���=�łM� L�@:����M��,/�X>O��a{�5�]�1�����7 ��7Y3�mHE������g5�麎��A��O�"""���0t��9��u��!��`��EA"���i�V+CNI���>b��ǩ��(��`0���T�:�ðlz��|h4h4�6%��v������� UU��fmL���I���N&I��6j���Ɉ�>M����[n��[�� �5��,�bH���ӦHDDDNp'""��������Y��<z�a���d�1���Á��)Ӛ^��&j�y�^$	Ӛ^�����6%���L�[��㣁&��h�|����s�� `3�S$fff����Y7��������6��I�~�%�2�N��,���������e���@�T�{DQ�����W�pp�S�n�����^�kY�������ׇ����RѲnqq	����tzz�N�mZ��!4]�K�����������@�`���
��>(EQ��xMk4M��l�CDDD�� ""�{����n���~����)�R�����́DC0>��l�;??C��i�v��_ `~�����Ghе�\������p:�X_9P�Q�Tě7����Dɲ����B����L&���C�5�D4|� @��_
$���S�����A��� �p8E�m3�$9`�>����z0�փ��4��C�u�z]�z4��^������v���:D4Z�v�_�Tjsss�����|>?��vP�s��ST�ױ�����W��/B�0��W��͞M�hp����׿�
�$���$	��+������#�i����WM�����7_������vqqq��陾5��"��@�{V*�JM� ɀB���Z��u]ʲ�G�n��6�"""z���NDDd#M������D.W��w�����RLt�n��O��t�]�l�Y,6�@�|�T�Q����M���DQ���e�B�����M��sɲ����&u�j5���@�u��݂�VVV?kj{�����>����p��ZQ8�N(�
UU?���f�����L�n/��Ҝ���;�tn���v�n����j�����3"���T*�����r�=n�_~�k���U�V���������eccq4�M�{wjS:T��������M�� &&&?lr�Q�d2H&S}k�^/����9|�.�H�&>���)SSӸ�����8�}�4�R	���ox���.//L���w����"""z���NDDd#]�����Y��<z�VWW���A��R�e�f�����Jk#Q��Ŝe���1'�����,�^���S���\�@�������և��&��_s��599������5�E��A��b2��A��
����	��Uu��T?6�s��}j�7�u�v�{_-�Z-�ZM4�M��m��$����
������G29>�������%n�y��6?���[�ǜ��A���u��n["�4����E�X@��,�۷G���_�l���d�Y~��I����Ź�=0EQ0>>���s�=}�B���$	>��J�o�����HDDD�܉��l"����v�v�J���	���ɻ�NL%�g�Lo���ʩrv������4���r(6%����������T*ِ�>����U�	ow��6���C�ӱ!�I�e���"���a8;{�w�ށ��'\.�n\.\.�ǆvUu~��(��{��0>6��Z-4����F�f���D�4��(X\\�$��!O���coo�z}�)�n�\�X^^����_@��F.��@��������hA����o���ׯG�Z�"�� O���eSS�89�X�\\\|���uqrr
WW���!�G�Z�v���:ʣ
���ݪ����v���1ѳe�;�����(��L����]&'�0==cc�������mN�$�O��D��5��'���~�����5�)���cww�����(:�����j����=�R�皟_��� �n�_�f�iC*�S0���lb���lbk�5nn2CLF��I��׋P(���8��'0;;���y�RC(�����$�ln!A �2\.|>߇�m�����16G(����8I_�56 ��h4��� �P$�2�����%����5�ny�RD"Q��}`�@�ZA"�0}�"�
A@�T�1}_�ZE29nzM�����&�kj61�  
��q8�v��V+6&#z�n?��F�QPU���oAR���s�R=_lp'""��lƟ�{5���+��~#=^�|o�vG��IE��kp8�D�t����ɍ6ZXX��g~������M������GLk4M���kt��a�z�P�5looq���L�cuu�4���\.���-�Z�!&#z\EE0B<��x
33����C29�h4�@�vک,���1�k~w�=��FcH&�155�����|>߇C��ި#=�^�t�(�-��|��AUU
����T*eȲlyXED�1�rY�z����t:�ayP!�T*rHˈh�A�o����u5�j5$�I�k�������4���n����� A��լ�0R �ľTDDD�܉��l I���������(�ꫯ ����'{{;��Gtϒ�q����֜���R����|>,,, �ѹ��`oo�S3G$baaf� pj���aq��94o��X���������%LO�|��0��������{��>��H��㘞������	��`��C�3o�?�.�~��h��)LN�n����P����<�G�Y�XD�^C81�&�}>��`�B��9!٩P(�������9����d���T*p:]&U� ���1"�j�x��0���F�RA��Mmv0�����H��V��D�H�����Ț(�Vׁ�,���ڮLDDD�܉��l ��_��w����&&���hi�����Gt�A��\��tpp���vZ]]���4�y����F��p`cc�,����9���ؔ�>G ����@�����dlHEvQU/_n"��=�v��ۜ�Gϊ �x<�D"H&�133�������D�������͚���^O��i�v;��z��j��n������0����A���<Q���CLNN!����B�'����h4������\�t:16G�\F��)�OI>�C0���/�2� nnnxM�)��H$���dY�$98�eD�@��A,f>�������ʦTT��1>>n1�݃��KS=}�a�n��OEE>�3=`(�┮�ac,""�gi���DDD�s�4M�7+����)��wyy�N�3�DOJ<����z~~�ia6�����k���M�������r�Mj��Rzxx`S"�n���5d���7U��`0��յӥ��簿��^�Ӈ�i�$	�@ ~ �@ ^�ϴ��3�N�n�N���fsM�>�����4�n@�z0�CS��H�A�pHE��×I��r
���    IDAT8���K�ȲE��68Q������?�3M�P�VQ��Q.�Q����ߜh�Z�^��/^�!���{TUūW_��������]t]���6^��n�۴���cuu��;lr@��6޾=��Ҳi]*�B.��f��foP.��ָ�$����o]�pyy���پ5.��h�̉�Q�\��i��3�]A@0D.��[�i�&n{�����h���NDD4d����N��X6UU1���Q{w�)�D�ILN�o��v��bd#Q1;�²���#���P(�drܲ��萇� EQ����tkŝL&�w�NmHEvI&Ǳ��8��d�0pv��޽�߹���\����~ ��ß*~װ�n��nw���NO�v;�~�����e�v�I��(��_
E��:����*I�gF��p "�k:3P�7P.�>6��Z��f$�o������R	KK��/EKK����8::�g�'���bgg_|����H$�/����M�h��5"��јI����e|���i���St||�_���0{�;;;�l���'��]^^`bb��5pzz��D��0�ED��o3|�B��i��aY���n���6�"""zv��NDD4d���{f�OM�<�����j�������S4��vqqM�lJDSS�PU���l�RɦD�}�$YNg���ބ{�DQ������
�v�<'�?�KK˖�鿯�ncoo�Jy�Ɉ��r��>4��(�o2�S��F��B��D����������,�Cw魈����w��	������	EQmHkE�������x
�퟇r��b��R��V�9�D�#�ˢ^�auu^�w��I&��v�����ôOD�����67����:11�f��)�������!�Ӊ��9~���-��D�o�$ɘ���!��z=\]]bjj�o���E$E>߿���>O��g���</E1}�m���DDDC�w""��
�>cV0mr�~���	'Tݳ�)�����S���r����89�ͶQ��_���7u:ڔ�>���
|>�e]�^���(��Ӆ��ux<�5����v9��=UU?4��6�r��.�v�F�f��_�h�n����w8t]G�y�����������t��v��r��v[��&UU16������V��R��R��b��N�=�lD�T��ķ�����>���嗿���6������*��v���a9e~~�f�bѦtd������kk�u��8r�
��M���NOO���$I�&p}}�F��+����8G*5a��LMM������u��-�;t+���4m�
�J�����| �"���=M��f���n7���WvFzԾ���\MNt�"�&&̛�/.�y��F��|�5��g��6%��]	�²n�j56�<433�H�R�u�v�_���'��`ssN�k�ﹾ�7{�^B����@8���$���1;��h^��d���0�l6Q*����p}}����x����g�d�(�V+h6��v�<�<B�a����l�Z��P�#�I�����r(��h4�v��$پ�N�$x�>D�1LNNbl,��A�=h�?C����\.�N��p82�ϔ$I��h�Z���6��ak6��t:�Ḑ�
��H$�\.�^��Y�F��q��P(�t:��|#�i�@(�[#TU�F>��EQ���D��*��2�ݣ��Sd��pX�dY.��[�2=7��NDD4D����f�OO�ؔ��+��(�J��A��LN�o��u6�!�ǃx�|b_����ٙM���dY���e]:}�P,66��.M�a{{�6��<ccq,--CŁ�u]���������/�ӅP(�H$�P(4����i=�ju4u��u�jU�j5y"4��j��j��."�n�^|>�n�^/dY�-��};e~|<�0P�T���P*9ݚ������kPŲ^E��������� w<v��Wp:�����)I��7��ߠ��ٔ��"���*�����y�gc2�sqq�dr.W���h�@ �r��d�������!�?�LOO�T��
��R(�H$G�Q�x<P�N�o�a�!�h_*""���DDD��u}Ҭ`j��f}rzz2�DOJ0B 0����F����ݯ/� �O�;9yM���QXXX�l2i��x��ئD4(�χ��e�:�б���z�fC*�����:L�n�����FHzDсp8�p8�P(������n�j�j�c#;�*>O���^�=Ԑ�|: �t:��z?4�����liz�@��g�V��B!�b��B�]�z����꯾����D��������>��?��'PU�x´��vc}}�_��ap�C��vqx������uccq�r9N	��qr�kk�u/^���o��)���n��Ng�L�o�C���Tx��>t:�j5x��QGy��nn2}�4m�@ӶPDDDψc�����*Y��DӴ���>�/7_����u���o9���-..�N+2o��q�M�� fg_��T�Uٔ��/�affֲnoo�F݆D4(Uubs�H�uC����r9R�09���c|||��)�J��z�f�����eccc��������|>$i��K4��J��l6���������	nn2(�Jh4|�HM��C��@�T��M��g�d2�T�h���u�,}�$I����crr~��������0i����TU����{<"�
�<��=�B�`�����,�(�6%#+�fN�˲i0"�N�h���ϗ����kh46&{���:R����E�qs�C!D�E�@ 8����!!�7�f,H�T�u���+�s�w""�!�2�逸��E��q;#=Z��8=�w�������y3u:���F���5��jZsp���/�v����e���%.//lJE�E^�܄��=;{��>����x�r�`h�ﹼ������Ar:]����}���D�1��n�Ə���tP(�q}}�w�Nq||�L&�b��F��fv��n���(�d�8??C6{�J��n��C�,�o��%A���F4���$"�(TUE��A��ڿ���0�|�N�px����r{�\.���6������Fc��/|>?z��ՊM��J�TB<7���p8�(
Y�H�QG2i~(������ʦD�[�׃�����`���F>����=�t:��Ɔ~}�)�e�b��ڡ(����6�"""z6��NDD4^�w��n�}��_���������^�R�M�����h��y;�}��K6���011iZS(����{���-,,"4�f�j�����0lJE����!�nt��8<<�!�����+�\���ɨ��opqq>�dD����bbb����E8����Mg�0P�א�fqqq��o����)��,��
Hh��.����<��.�N_�Z���iCEȲ<�?�TUE0D*5���1(��n��fwzPj�*J�2���[z����8�'?r���X, OXn��¨ժ�H�@��Z��D"aZ��zQ�V���@�Ӂ�����[#�2��j���ɞ�F��Tj@��}�,!�����	3N��t�/}���P��=0#���DDD���DDDC`�?�u�7������ش3ң��v��~ϦA�{�v{0??����������	������l��v�`6�`��UvwwxC��y�b�dҲ�V�agg�������Xkk떛��mlm}�R�8�dD��x<H�&������A�i��D��D6������qyy�B��F��m4r���^��P(���
�(���t:E�r���%�
�� ��SH$�PU�6'����n���f��(�[DQ��X�a�\.ې������X���� �D"������@�Z-(����W @ D:}�k�#P�V�J�L�|��)�|~��������eq�ݸ��A���sD��0t�B�Q�x$IB>o�uEP��iڿ�+�s�w""�!��������"�񸝑�w����It���L׽��7{�!j�Tj��� ����+��&�lllZ6^\\pe��'077oY��t�����}��MNNaqqi�龕J[[��P
����D<��0�����5��5�_^^����߿G>�G�Q���=l�a��j�X,���
WW�&�w �P�%IB @*��8ٽ�a�;����ps����1m��D@(���B��z>�f�	M��7����p8���_��r��Xl��=�$Ip8(
6&#�v�,+���Bp8$h���B6i6���� p8VM�D4�N��H$:Ж��N�e�JEӭǂ L���6�"""z�N����y<�D�����j~����t:���}��7h�룎A�$�\.,,�7��9\^^ؘ��r8X]]7��l:vwwM/��p�x1�H$bZ�j�����I^����ںe������z�F�aS2�o� `aaSS�O6{���m�N��Q��8�������P�s5MC�P�������w����k��N����h4>Mx�d�h6�0��B�{���MvO�&���p8�j���D#a����`08��x�^���r9n-z�*�
TU���w�
��fi�χ���M�Ȍa��kH$̷���>�E��m��ѝj����q��~�����u��[��A ����[��x�ɤ����Ȳl9�n�z=�j�����g �����������������������˗�v�y��:����F���x�b�r5����P����e���9�����׋��e�&齽]6H? �����WM@���b����B�������<�B�E�h/^�aaa�p�������j"���ݻ��&�Z���z�z���*������X,���B�{?@�(
��0&''
�!��_[�v�R	�f�Hd�-6.��H�|��3�B��@  ���' 8�.8~�y Z��N'�^��	��&j��)v�u� "��E� �g�&�v��P� �[��I��!��:ƣ I2r��Y��(JSӴiW&""���DDD�L��0�o����񄝑���Cd2�Q� zdY������b�����6�z�dY���鄨^��7ov�Z�f� `c�eCT&���ŹM�����6�ġw�NquuiC*����N-�u��o��J6
�033�����q������)�GG�x��=
�Z��m�Yk��(����B:}�F�A���{��t:�D�JM��rC�4�Z<(L����(�J�F#�[��(��h4��=N�|�X��P��@��2�2J�)�K���$�o��(0�r��d �Z�D��w��f��A��B(6݀��xpuu�k�D����"��F�-I�P*M_AH���m�EDD�������~� �	��wM��L/��'_�{N�&�'��S�¦5��h�Z6%z����Lk޽;E�X�)ݙ���<���v����i����јe]6�����h\.67�������ickk����6N��X^^A*5��kz��s�z]d�Y������2�4j�*����ij�*nn2���@�V��p:U����E^��D�d�$��j��l�n���f
��"I��*�
�m~��t]G�X@<��|�GP,��tlJG�躎v��Xl̴. �����À��[A�,[N�{��tL7����^��J�lc*��K�$�M#t��� 4#���DDD���DDD�HQ���i��������˗�vFz�
��vwF��IE������*�
޽;�1���r���d>M��nc�'����rcuu�r����>�ժM��J<����˺j����m�\=R�@ ���,�+ܩV�x��;4��!'��N�b1��-`aa��'��Z-���8==���r�,��}&�0�h4��eqqq�R�M�AQ�{���$	�`��0�f ^ixz�2��^/\.�e�(����l�Ѩې��[��E�V��X���� �¸���p��h4��z�v�?�+|>�in4�[�VC,6f����P��Ј��&�ј��-�ۃ��S=]�n��ݒ$	�\άD�e����o��DDD�Ա�����~���a�=8��`9�n��C>oz����H$16�� �}{�F�M�vX\\��>���1�ՊM����ښeSH����)�<~�kk떇��6^����T�h4���8�5 ��9loo����C�˅��i,/� �H��r�d��gi���d�899�۷�(ܲCt�Z�
�.//��e��v���ic���\.�bcH�&�r��j�8����0td�7�e>�߲��p�A@�T�!!ݷV��^��p���i�n"�7776%#3�r	����}UU��vx�~�ݎe����B&�v�u�tS�$Ih6����OR&��h���Y����I��b�M��Y�q]���������46��/��&]_���Ȍa���~�&4�{���jڨ�j�ptthc�����c~~޴��h�����Dtg|<�Tj´F�z��ނ�i6�"3�����W��h��c{{����Tj�����M �wuu���}�T���k\XX���<��醜��n��N_���ۦ�B��v�}/��Dd���T*����c���:�e��(���|O!
A�u4Mp�;C���a�B��AH��b�0�d4�jN�^�ϴ��rAE�E��Q?�����!����Ad2i^{�Y��@8��:��8�.T*�ZM�=O�F�D��������ե����.Qt��>(I@��5=\cF����I""�{�w""�{�(��iڿ��q�χ��WvFz�2�4���F��I�D"�M��ޝ�R�p;�����4?�tp��i�6Skk�SԀ�����A���^�ײ��� �|ކTt�&'�077�A�b��''o���%EQ011���U$I8���^>G���AS{�Ȧv�Qk��(���@�T��ip���r���t"C29I��h4ټH��\.�Ѩ#�Zn9 �? ���-��T�X@8����u�@ �F�Fݦd�O�VE 4�#�"�n7nn26&# h6�H$��5n���W6%z�A@(����(�?{wٶ�	����p4��q��3ݧ�9��B�����J�W0)	$x��f� !��PT�*�B!�jX�to����v�v8"���{3��{�97c�p������^q�_�tD쵿�}(�vEt����'����l��v6Y�֤�i��DDD��������(�򗚦u�;5��X��H}kue��D��ٳaV�����:t�{���a||B��P�����A�諙�Yi׻B���m��/���"�.�y��n�����ƻZ��67בL�6=:���������|�nΚ����������y�E�D�T�����e�{�p���o�l6cpp����x�h��,̢[U�VQ,
����:0����A6���@��u���Fc҃8�@�\�Vˠt�I�XD<�:�.J��F�.����ݎJ����T*~�Y�V!�����vK������yNxX�d2%4M�Kc=X,p'""�]��[�K�|�Ng�Q��i*����4Nn#�)�ۃ�	qA�����9��33sҎ���k,r3X ��'�MӰ���V�iP*�F������+�X__c�N�Q�ӳH$��Z��*VWW�Ͳ�(��ɄX,��������v�B3`ss��	����L�^G6�E*�D�V��b��4EQ�r���G��:��*�Э���8?�!�b��r�\D6��\�Q�6J��Ѩ�7��dB ��Y���k�/��~�:�o��'|�V.��H	���H��Ž�t]��f������t!�����-P>��]���fS����z�i\"""����DDD��b������k���ŋWFF�[�d��w��A��������u]ױ��&�4A���H;g�� \>�_XX��j�;8�G6�1(���n,,,BQĝ(��&>��v�mP2�&��������ɟ?D�P�q2z�VFGG1;;�H$��v��f�V���677�L�\.C�Y�D��4MC�\F:}�t��vv�C�{R�f�!!�H�l6�Z���A�P    IDAT>�n��j���~���5�Á@ �S�;����z�M�����,�n7���JF��E�A�l�;��f�L&��lLa�V���!��g��P�Vxh� �jCC��<���T��D8��C���l��yN��d�ٶUU]6*�C�w""�[`2��RӴ��8���FF�[+��,R"�v�Ϟ�7#���H�OL�x���I�{�X[[e�!����#
�T*ll���D,+��^�j�躆��ϨT����X,,..I�~U�T���G�jO7�t:1>���s���0�o�]�i��vw�����B� U�a����n�P�@2y��ↁ�� ���l��� ����t�P��x�@7��*���p��]M������8?��h�)����p��鄮�(.JF��JE��	�ޝ��E.�E�ɉrF*��]tq`w��m�g��5���$�!]��t:�p8�:ʽg�ِˉ')��4�10у�w""��3��t|����K���ܬ����q�*�-�����\�2�A���
ל�����N'fg�$it��,��h��:������jgg�����f���/�z����˟�j�;�����arr
O�>���q��j����/��XG:}�z�~KI��4�M�r9�RI��u��M�Pn����� Z�uѵ麎L&��)�����bE(tY���%��I����� ���ܱf�	�����q����S6�0���a����t�G�Zm�ժ<\o�z�.l �(
4M���ݔ�����]��D���M����¸DDDD܉��n�j������f��v��^Ǒn]8:��/��w����f����d��90�?��ё��/Y�v]ױ����F�����%>|�J�pr����(�������S�����n�����R��As�VW�ٙ��IA8���FG�000p��4MӐN�b{{���(<�K��i��r������<p�n����p �"
CU��"
��td�X,x���i��X,�Fc(
<��Gt]G>�h4&�J�����,���w�P("��b�t\c�;�h�Q.�LF�r	CC����ۍT*i`�ǩ�l����pt\�v �JB�u�=<�f�pD�l�.)�	���h��n�PUuӨLDDD܉��n�d2�#Mӆ:]��ayA˟?�T*�u��744�P($\����Z�fP��+
cxxD�&�>���A� ��0FGǅkZ���VX�xx�^���J�P��2VW��0���\.�x�R������S����=�+S�hss�H$�n�U ���|���~vv��?"��F��\.����N�V����=�͆p8�h4 �T��N�+��ϡ(
�� �d2!���w�i��(�ˈD��{(���ǋ�������t]G��@$�����{RU6�M8i�j��V��R��^k�[�D���Lf4>_"��N��c�{6��\V�ݬ(JHӴ���XDDD܉��n��u��w���%x<#���f���?���Y�R��s��O�J��;�z�fg�Et��cmm�v��T���d��¢�o�<R,JE�X�V,-���".k��������������K�l�'\�\2y���- ��H�S��(����oTX
���/������-
��ND����=�J�X���d�����&HX,A�b1�����R�*...�j� ��~-r/�J��yH�_��5���/\�����Ņ���j�
�����q��d��bA.�30��e	'����R)�^����"�����r!�dG}���������(���FR1]��+�2=D,p'""����7�����t�b����(�.����c��H$�x<!\���Ǳ��#O�8==A:}jP"�'O&�k
�vv�JD�)��_��u+++��G�n�O���u�>:�Yt%f��������nT��n��N�bcc��G�V+�����z��L&�t:]��r�`6_�1��B�D"�ٌr�̃7ԵR��Z��P($=l�(&��T*�jU��M
x�^8�����������J�"������q#��sz��TU��b�����b��^�s�� �==�ՊJ��j��UD7�l6��l��� ��w����j��������5������E�5M��t}xdcc�&�_?}@���D7�������p��&��6�����ɺ�k��n������
뺎��e4�M�ѷ���!������#n�ϟ���xww���E��l���(���
�a6��u��j5�css�l�V���c�n����L&�l6�r��}�l6cpp�D&�	�r��{ԕJ��r��P(�E���p8�J����>r~�C$�L0S�N�AUUò�/��m(���AQ�}^�'')�r�e�DbHX���J����c�J���:���8=��M9�!9l6;2�����l6�5M���EDD��������f�g]�;V/�/,��42O_j4x��ǻ�A��|�A顚/_9z� �h�ĐpM*���ٙA� ����t:�k��cK������F ���<��6JE7��x����U�������i�;���tٱ}nn�P&���<K��������R��""�)]�Q*��L&Q.�`�ڤ�W;1���#�,�*���uvt'�Z��B��PHޥ��=�j�E��B�4�E�b1ὕ�l�����Y��t�k�R�pDx�d���j�P*L��i���,|�c�X�l6Q*�L������}�8���t@tC��#�u�{OQ�jU�$������Q�����]��j]RU��;]7�L����t�Qӏ���R)Ng#����)�\�k����u���1EQ0;;/| �i��W��@�h��#�5�fkk���cV�KKK�.�����ϟ�w�'|>�?_��"/n�4��+�d2$�~�(&��q,,, �;�����α�����}T*�,EDƫժH�O���`6�000 =��-_����I8��N2�F�|�pH�]�(
B�0��:�/�D�ـ�j�"5��EQpq�7(�����j�Fc�u>���i��\.u��=����V����f��@t�V���ty�P��TJ�u������v�``,""��wDDD�d6��;M�;]�'x21id�����{T*���A���v;�>�n��X� �X�x\�&�<�{a �ق��Ei�����evۺ[
�v{��t]���
?���A,..�lZ  UU�����5$�(&$	��/ �v�o�[4MC*����R�$��ѽ�l6��f�N�BQ��P�����f���bqh��r��Ew�m�f�\�PXz�TQ�!���b���-l� \N�JE�j5��ѯ��5�10���2�L��m,�5��.���f������*�N�p���r��䄇@�n�n���r�u�{�f�"�O�UŬi��cP$""���DDD���u]��<;;?ǷI��u���c����1�C@�����a�#EQ0??/�P��*��lrr~�_�&�?����A�����'���D ��`�����������v�˟Q,��u� �b~~�hTZ�׉��q||���5d��>"�{��n���'''�un��Z-�� b�Z�6RG�V�l��"�P(�S1'	��|�������@ ��3v�K�b�xB��?0�F�P@�^70��V.��H$`2u��u�=H�R���c��e�NE����D$�i��]Ǹ�L&��2��f�5���u]�c=,p'""���o6��I�늢��~8ҥ��=�Rɻ�A��L&fff�Ń�\�k���Q���1�٬A������p���kXYYF��20���7(}� ��<���m�R�M��,.v_����'v����~?���H]����j�Tؾ���4��[Dt�i����<��$��&�nOW߭�f�X
��D�j�P��Н�X��F.��� �� ��&'a�M�P,�Ƅ�\f���t��t�s��B�u����9^�'')�R��iPE�@�l6��n�X�}m/�Z-�|>8�Ύk�N��cS=<�f�`�Z������=M/�� G]�]��iڿ��b(Ƴg3F��[�>~`�0��D"Ңꝝm��1�K��`nnAX��*��V�i������9�(�/_��p��]�X,x�|	V��p`�����'����w���,n�N<fg�06�6��Z��f�������9����/麎R������&��:�c�ZGP�U�h�Ƃ~��n#�� I�@0b�{�h6PUUڍ��p@�4
��tWJ�"�������jC�����e��q�}���F*�d�k�UD"ю�-*�2�ժ��������0s���jE&s&Z�X,���i�ܨLDDD܉���AQ����`��O�N#�/��u����c��g�f`��;^��j��e��^�Fc����5GG_p~�3(�!����4u��������������u++��p�x�><��Uq{��ħOYE��t�ٳiLM=��ѹ3�H�����67ב���,l'�����=�����z��v��X(��h��=HK�JUUd2g�]0���klb�J�"��"�?�!�;T�V��L>���'<�i�˽#E�]�l6���j�b���7��jC:}j`*��GU5��qt��_(\�L&STӴd`,""��t������KӴ1т��!�����#ݐ������8V#(�h��8>�{aE1arrJ�n{{��n�w)�#�H����`�Jq{���ǏQ��HF��b�bj�)�����>���lbggo���T�?D� i��T*�7o~���m4��k�w�����7��z�U�nz<��&>��eѺ����kw��67ץ�E���\W��7
���8�b�J����z�Ldtt��2��ґJ%�+��y�H�R)��j�u����u� PUulBKDDte��$""�"���4M�띮��n,>_22R����;;�Г'p�=������uv�X8��аp͗/����JD###�D���|{%�oq:]XXX��$~��e���I�������/��"�l^vn�V�[�.)��x<���E��(ʕ��V��GX__E�P�aZ"z~�ѽ�h���^� UQx�^��	 ���,?C�rO��,�? �\�;
�¨V���w�麎b��X,&��e�Za�ِ�eLG?W(�'�����l���z�t��n�XP��Q.�0w/U�Kp�&����v�\<,"c6�e��LV�uOӴOFe"""zX�NDDtE&���4��lЉ�I���ѡ4����c�5�ł���&���	�ٌ�����9��~UU���ƃ�Zm���> �u���| |�E���s8�N�f����������n7��^�b�w~m4���j5q�Hz<�XXXD<�V�PUU�Lcmm���,l'�GI�u��%����l6��x���j2����DP��Q��z�����i�d�����.r/����w�5�Mh�&,� �ۃZ��&%wD�.'�����'EQ�t������T*��	��������8݌�ip:���/.� �zݐ���w�޳Z�8?�	�ŚL&��i�ԸTDDD��������HӴ�����/]::�������$.X������x:?H.�R�ɓ'�ҩT���ؓ'�z��U:66���s��Թ�����߳`�  N��XZzq����˗C����{{�h��=HID�_�����~���a�E'�Sv�ca�9\.WRR�i�������t��(����N��;>>ꪳ�ӧ�p8$�o9>>��?��~��w����D(6(��%{�f3�јAi��J����.�|>�uMӾ7(
у�w""�+���]�4[��6��07-�q���]G �s
�!ኋ��`ttLx]�4���n7b1�$�v����c�7bxxD�����|ހDt].�ϟ���*/no6����#�����>3�-��������`0t��뺎��~���a�Z���AU�88�Ǜ7�E*��V��`0�����S�����m|����"w�Ʉ��E�HF7����f�)\s9Ap����~N�5���J�MM=Ny�ەLK�Cd{�ts�r�bQ�fhh ?���K�u
������A�uM�\V��;��=W��KDD�)����=�t}dd##�FF�K�F���x�1��Z0�����Z�H�^��ظpM*�D&�1&affN�S�foo%�_�X,x�|I��\.a}} '��WN�/^��������5�M|���K�`0������*����X]]���ɵ�=6����<���3�l�+O�P^��D�v���fz�4MC6�A ��T�p�B�8�W���Z�"�
�9h���;R�V�����V��v[Z�K�C�4X,�|��m6��'����k�n�V��b�:������s:���fC6�.6��NM��c�5�&""�M�����e'�9>:�V�0"�Yq{��@6�5(��%�Ĥ�:��(��w�V�H��%�oy�lv�x����X__��k������x�|����V��ϟ?����s:�X\\���"�v��__,���|���J�	���Z����U���Z�=-+�=�Ƌ/�\$OK��§OQ��'ƙ�f,..��������<��}���x�>ѷ���H����ƻ��E����Hz�vttܘ0���YF:�bhH��NDb�R�M��(
<�p��i��Aq����u��p�i�ֱ��dB,72R�b�'��8�N�"�T*Ń$=�v��]K��S���TgE1�ɓI���m�mܡx<�p8"]����b�{�j����p8� ��ncy�*y=L&�O�L���@ p�n_�Z������
N� "��R��O�>`ee���o�|�x��{LLL�l��Ǫ�j�T�.�7d6[�����e@2����]�EQ033˿�;R�Tpzz"\c�X0>�ĠD�j�������x�nF�5����� �o�u�"��t������/""�.������K���G��h��Q��j��N��u��vٽ]�x]�u���7������u]�������ȈpT7 �r9�����~��pbrrJ�.��HL�ݹ���]�R����ϟP*�HF�Q0�������1(�ն!UU���޾}é4DD=��e��o����v�}��*����Q���o��z���f��ϟ?vu��*$�nh����Uh�x�����}������pM<����۠Dtt�E:}N6�n.�LJZ(҉�D$v�)P�Q7�nl6��7 
у�w""�.i��7Eׇ�9֕T*)}PBD��Lf�b�i���͆A�'�˅P((\��f؁� 6�M��P�u����������i��F����M�2�U)�	���x<ҵ�zٹ�T*����Á���XXX�F!�����y�[��ށ���t]G2y�7o~����O��옙�����aSz��>~��U���n���/`��HF�Q�T���']�'��D�7���kE�!5����k�~W�t}�fCz0:O�d�
��*��ܣ��b����p��ibP""���w""���4MV��Y�ޕ㣣��@�ע�(,�pM2�4(��566Q} ���ۍ2>�DZ8�L�����7(Y�ccc]ڍ�(��������4++�(Y����	|���^�T,���{lnn��l� }K�����&޾}s��G�@ ��FFF�(��$zx�:>���A{�Ӊ��%�ݝ��#���릧�a�p��]H&����ߏ`0dP":::�5(��J���-"��Ai�MӸ��%١&UUg!{�DDDD X�NDD��������{�������OMSqrzr�1���А�0M�\F�X0(���p8���r9��%�=n.�K:ՠ�g�;.���O��|�������:��g���4M���2�?B.�/_�³g��CG��hԱ�����a)��V�X^������+��d2abb/_��� ���Z��O�>�ՒVu�ݘ�_���G���Ɔ���͌?�    IDATf���S�����Մ���I:2H�VC&s&\��v˧���]\�Q�T�k���JC�0
ܻ���^�u�l����Aq����w���������]O�FE�k''�hw񠋈����IR�c��<^���GG,�6ʓ'������
~GE��̜�x�T*��`ߠTtU��S�Fc�u��ccc�EQ022�ׯ��v��5]בL���HB���8�l?�����4�J��x�x��;LLL�����V����#��t��ss�,���Z�&��6���(B!�!X�}�\N:q��ruuG�㲱���������������#.<%��
���#���U<�FӴ?5(Q_��"Q4M{!��H�;*ӥ�㣻�@��b1�a�v���3����n�>��ȣP`}#x�>�B�ەJ'')�ѯ�����w(�4���q�t7���1<<��ڭ�Md2�'����v�ի��*b,.��ݏ��ن��=JHDDץi����i�}=���w?`p�ߣ�t��e��.wU��0==c@*��\.���S�gϦa��HD����#����F�V+�fs�5�pN�ˠD�S:}*=h��'AQg��rrm�dM 4M�+E!""�k��%""��Z���4�.��P��jdt]G*���D�e�X�|֜���@�ǆ����|a�v�LLLJ����p����n���I����IGH�݈����������8�&�	��Sx��;���C,��l6�����?�o����j5,/���*�ƕ^�t:�����O��l6�(!�7X__��>,�uu_Gwcww�F]��j����i���U���v����ts�=��`|?zIUU����9�H��K�n��}��E���n�?5(Q�b�;���]����҅��ٕ��t��.�J7c6�����JE��y�=n�P>�x��������Y�&�	33�P�o�B��$��K�`O�>�j���'�<"��_���(�r�W�H�O������{����z#�9Û7����t]ޝ�$C?us�Y>�_��,67�ȋ�GFF144��Pte�v���u�P�HԀD�k�f##��Z�%zܺ��Fc�z�c������lF81(�����x<i���ifP""���j<"""	M����DB\�H�X�Dt3��xt��E�Z͠4�S<���b�9<d�v#(����	���]�з���c`�-\��*67��a��x<����x9�J��`߀Tt�ń'O&���+�\�+��\.�ݻ���XG���QB""�5MSqp��w�ޡT*^��KK/011�F�D:����NWk���
qB�}���j����3����R��ZM龻�b��|�ݎ/_��M&����L�ZA�(.����{�D�Y���D�.�L&����qM���Aq����w����\���Db܌���1��]����G����Ġ4���(Ҏr�j�\֠D�[,����pM&s�b�jE7t;�^/FFF��vwwx0�r8XXx�ո4���HEwm`` �^����ؕ��k�������r��	���H�J�߿��֦�s�/)��������,���1�|�� ����9x��)]t7vww��n���3%��;:��f�)\344��iP�����B��H�W���ʽ^�to��:+.�:B_����4m�|��������j�t]�X��1܅��sT�<�Ot]�I�v�,�{)
��p�qR�L&�ƞ�躎��=��ϙL&LO�H`��<NN�#��xV���K]�K��ϱ����2E�Z���n�a�_+
x��G�C׵%$"�����$��o� �?��+].^�|���I(
S=t��{H&�/L&�<)�zO�Tllȧo���B�}�����@�FQ�{)t{d]�m6�ѨAi���4��p?���O6%�.�
�u]7�l��kP""��ĝC"""]��-��xbȨ(}-��C,"�6�ɄHD��#�>��]�k]�����z����Yڠ4�����t�y*�dg�;���\.q�v����u�Q��RPT(���Mc��C�t^����nckk?�G�Z�aB""���:>����u�ۭ�_��իW��A����A&s&]g�Z���V���%�X,tuParrJz�N���$%���F�|h��'��H����Gt?��F�4��N4c'}�k���h4�w�޳�l��ō�4M�w�ICDDԟ�����H@Ӵ%�uYWe����"��p8��"\sz*�J7�����z�k��$=`�X022*\��*�|94(������аt���6����{
fg�]� �V�auu���h4�ׯ���#����\.��o�pB�#�N��͛7H�O��:�ۍW����w$�3������ҕN����a6��EW����JE<��b����i��W����@6�N��Ą!y;]ץ�D\.��A�'�}��jE02(��S(��{7dϖ4M��AQ����܉��:�Z��4M�x��n�#�/U���^ѷ���Q��b�r٠4��eG��4ME*�4(��666.=�qt��fӠD���(x�l�"�>��e�\�D�755�P(,]�j����	�V��Y��X,��-`ff�JEe�v��XY��,DD�X�����:VWW�ju���d2aj�)a�Z{��kX]]A�"���x<�����_��4M���:t]���#���2��Eq�����Ϣj#���H'����'F�͔J%�y<�&VD�U(\�u�� k�i���p<1(Q�a�;Qg.�������$�>����r���a���r:��ć�NOOY�i �ÁDbH���j���ȠD�s##�p���5�V[[�%�n���v�1UUU,/��Y�����������~���o����3��w""z<��~��2�̕^����?�����m��,�ٔ����zj@*��r���Դ�����t���d]܁��I |��k����D�o;8��������~?�N�Ai��J���"]p��0�ĥy����Aq����܉��:�4����Cw���Q�D�Y,&�ޮ�*��zlxx��~���t;�ǟH7����A��+�˅��q���-v׿gB�pW#�u]���J����h��`|�	^�x	��� �?��mlmmby����i�ZX[[����
_�V�cj���?��z��ϟ?��nK�&C?ݗ�}rxx(��o��099eP"��P�@.��q�݈D�a���1t]��M���I�O�i��h4fP��G69�.�U�3����CDD�w�;HDD�mMӄ����k��8;K�u���(&�b�ϙ��3����0]��b�~�g�YT�U�=^N��HT��V���$eP"�ϞMK��r�2ȹO�n7fff�M羝�md��އ"�9�N�|�
cc�W�N�����?�s����2�3�}�#�����644��/_��r�(ݥJ����i�' LNN"�����677��p],��0(}���#}o�ǟp:����9I$��n7(���n��Ɉ�3������P`�{7<�𺪪�BDD�܉����j��{��w������RIh��A��P(��&\szʢ�^��l�9>>2(�����������.ݾD"�oP�FU����4(u�f�aa��3 �J%HEF��x��;�C��SU��[���#�z��C�l6���[[W:��v����w�FŇ]�?]\䱱���J��s�y&�^�T�j�ݳg�]�w��V�H�O�k�N'�����(6(��$�C��lx��:���wA�����f������}������z,.l�N?I%YEt]���s�R��X,���1�LH$��kJ�
��=^���5�R�LƠD���fǓ'�u���h4$�n�L&��/v�!��,���}R��E���$��`�X�~]�T»woy��������o��x��(�ٌ��9����db��C���M�ٌ����F d���}�j5��Á��qc�����C�T��)N,�J��|>/\�H$`6woFWsqq!��)ۋ'�o�4�R�c�{�6�x/VӴנ8DDD}�w�DDDߠi���x<nT����:NN�]��:�v;�~�p��z+��f?8�u`��1>���{{{Ƅ�_x����8�P����=3==�Wޱ�����O�v^�x����+�.�<Ƈ�Q������d��:>}�����+M`�Fcx��5\.v�~h���p8��� ���6�MS��%��5<<��c@"���l )i>�p8����d �fߋ;==^���S"��b�p����+�-�i�_1(
Q_�.ѯ���IM�:>-�X,�BFF�K��3vk%��x<E�\Ыi���&z|��ţ���:�Yv�5�ۍPHܽ�P��Ņ�ݾH$*�=�iZW�d���qD"Q�J�����:G?$�`�}��^_ׯi6�X^����m�{ "�[��:����������?�r�ի׈D"=LGwagg[�� �^�=�6 u��"�t�T�FQLO�����}����k���yh� ��9T*������P:}*<X�(
]ܻ���h� 4&Q��+ѯh��g��h�#�����}�|3=�͠�j���	p�$��W�6H�sٽ]l_>Ξn��j���t���t4'
c||\���jauuYZA�CQ��?���,kׯ�f3x�����{�����b��w��^� ��l���<fffY���躎��i(p�����h��vvv�l6�k�|��j�p||,\c���'J��%��.�����z��l"��
�\Nn�!��j�Z�����#=�d�X�Ԡ8DDD}��DDD�����.����$#P���� �v�p�ɉx�*��А�{����cm��<�A�|��A����)�l6�r����/%"�ۍ��Y��꺎���+uR���f�ai�%�����zMS�������#"��S�6��װ��UU�~]4Ë�`��{�����m��,w��cbb����H�����t���8�N�����#����ˣ�cl�c�t:-="ۓ����;N���a)�w��3����J ��Y����	܉��~EUUaK�x,nT��U.�Q*q3��:�Qq��z�����n��Ӊ@  \�J������'�kؽ�h>�O�9��:��68������XXx�Y^������y(�^^��>����T*�{�''�&#""�c���x��G���_��x����,F{@����V���P033�[Z$D9;;C6+�l2�05�̠D �v�����6�������iHI���|��?�5����Ѩ�D�Q��=,�b�#���+��iڢAQ����܉��.% ���l��u]�tZ4�v����?�6j����fB��p����唎�nu]G2)�L7����r�;�LQ<}*/F8>>B�T2 �(������:�}������x/^����}W�t�>�C�ʱ�DDt7j�>|xw�{.�Պ��_`dd����HylmmJי�f��/�j�������%m
�JD��=�l2���XW���fR�$4M�2(�c�K�=��0']C�RA��)�2I���iEQ~�?�� �Ǩ=,p'"��*�O � � � �7 ���E�8��w��D�#�@�u�&<]��d�~�g�4�=^��O�kz�~axxD�I�^��G�>}�O����<���=Q��L&<{6�gϦ�(�m�i����mll�CU�'$""���������,EQ011���yh>��']tp8�����t>�N�i6]�WLM=�ߪ�TU�vq�Z�H$XX�k�V�tZ�&��b���^9=7��l@2(���f4rN�K�>{  ��� �)��������U �� "�G��DD�X���]����O�w���X�.�n��9;��D}I65�ϣ�dqu�t� )���^��|����5�l�7̍d��166.]�����{"��4�B�Z�`mm����z�n�ci�eW��W�j��_�S.���޿�J���k"�^�x����dd����r9�:����!i2F*�B�X�����nO2y�f�)\322
�Y\tG7�J��L&3b��Ai�z��B�B�F�GOD�����W�?��N��5���#�w""z�b�CA�*��P�>��E�񐊢 �ƖL:�fa�5��v�������K�SU�R�> ����5�{�n��Iy��t:����A�H����ٳi�V����e�jw�Q�������w�z�]���,����^�p����H���A,Y�՟s��x��5��@��t]���**��t������HN��֦� �儰�2���8:�"\c�Z1<<lP�ǫ\.�P�����"�c����l�!z8J�"ht����j �ѹ��5XHDD�܈�衈Ⲡ�x�_��u�0�L��@0�M�.���ݘ�:��D.TUE.�5.�#������n�{~�_z�#�9C��bL#����a�UmcooנD$b��07� �I��iVV�Q��JF��ű�������i�������ѽ�i677���.+��=�Պ���b�f�SU++�h�Zҵ��3,��'*��tEQ<}�̠D �T��x2���,vqﵔ����D  �nH�wv�a�+�PU�M���S�.�������p���/3""�W���������+��P�KbQ�����I�#�%٦y6�aZ�����m���J�x�����뺎��c����SSO������l��S�)����y��v�ڝ�-��qt���?�����-�f��O�>�7;��t�>�C�^�j��(��z�g�f�{~t���5���J;���f��/�8��88ؗS�|�,"5��i�.����#%z�2�3�J"�CZ���mi#�h��MD�!�PA��Id{�7����� �/����7FDD�wX�NDD�"�o�7d7*h�5�C�h��2��EWc���<��˘lt*]��jE($�N}zz�=688��'\�ɜ�Z����FG��r��k�咴�crrJ:��wrrb@"ꕯ\cc�]��P(�ݻ�(��FDD�C�r�߿E>��k��8��^�j��0�Z>�����t������<5���v5�krr��tr��<�{�c��K�Ƀ� �A��tZ�������+���ԍn��ߒ0��	�Qc�;�W�:a��G7\��G���B����|�RIv�$���dBD����ŅAi�DbH:�1���[����	�뺎��c���␑�Q�*��[���N��F14$��V,���c@"��ݎ/^]����$�O�>��l�0Q�Z-,/�v!�9�χ�/_Kn��vt��̙t����!@ꝳ�4���p��f���x��M���ˡp��bA<�0(��J%%{)
	��r~���������u�=u�����jn(�_��ಡ�? މ��b�;�n�����?�
�{��%+l��0�̽�� �Nؽ��EA8�I��,�EQ�����Q�UJ�8y<^���t:�j�&'�J#�����=�v{��ٌt]�����J/�P�y�>�z��nwW�5M�����6��|߉��a�u{{�X[[�zҖ��īW�{��ziss���ccc٬�>��ޔ�$C]����;99A�^���k6��f3�5�x��C��.=4�D9����]���H?_d��$
�O �.�3R�,x�S �F ""�a�;ݕ��� �a`A�UEc�� �j���f�:Q�����l�5���t}�Pv�]�&���^w	�u]�a�nW(���Z-�����:1�͘���>��ukk�h6������FcXZz!���U���Ǐ�qzz��dDDDw#�9Ç�P�պZo6[0?��Db��ɨWTU���g�Z-�J33�p8���j�����kE�ӧ�%"]�wq�Zm���%z�d{�����1
]�l��n���4(���f(rf�N�x�������� Xމ���WŃDD���sA���zw� �c�����	��]�l�i�\F�R6(��H���u���J�8�\.�B��z�L�]�d2�099%]������    IDAT��v[VXB�6==�K�@ vv�Q(\��zall33�]wo*x��-J�R��ݭJ�������"����B�g����q2�z����5�~��b���<��B���ၴc��������ٻs�ֲsm���(Τ�A�x��]@'v�7��9j�4p��С:��?1�m�#G����ֵk8��Y�Iq�aw�:�t���6u�7I����U���Z���t�����}�?&+����z�n�Z���"��D4�j�ʉ��B!��1�������EDD6�o�DDd?���ߢd�@�u��)��^��h�&S���!��t���;$g2i����ߏhT݅���d\6ﬕ�U �n$GG���B}KK�b����sv��H$�L&�i�}ou���Q.���_���K+#""�N�|�5NN��7KK�x����c4^J�"����u�P��0j�^;;[���8�N*"]�q|�~��z�H�RUd_������`�pĢj�G�{O$|]"P��e�&����6��x�������""�;�;wDD4,~ ?A?�~=����ѕ�&d%��Q��(i�p��H$�p�6�u�rY���R��c��dSS>$�Q˅B�;[���biiY�F�ulooZT}L(6�y�V�as�Ѱ9�N<}��������}�~�j\����L�������w�/)'	|���p�Ǧ����О��K�d�|>�B!�\��x��4<���h�՗b��Wx6b�t:�N��\��`�;!&�� ����Ӊ���I"�>N�A1�0�q���� �3��w~�#"���wC""[>|?��w �C?��]iÕ��BI�RA����D��F��%�Z-�����%����,��E����xPzx���VZ[[;S�������r�\x��x��n����7;O �ǃ�>�ffԓ^��v�x�ꥡN�DDDw���)���1,�^8���H�`D��ݻ�h4�aj�gAE����%~712Q�����]�}>/������"��m��vqq���s�i����RQ�]Qjc0�L�u ?G?�~�~��� ~`i�u�c�����r�w0�.uu���(}��ID���N!U���7��R���==5>ޞ��x��r���p��a�w�n_��`ߚ��>|d �����׼(5�|>>��G�wy���_��|��ʈ��&C�T�?��_h6��3 ����G_ 4��K����������u.�O�>��.�w�����ԗ���IU4'''Ⅰ��U ��(''�Pu�4C�&���c�/��l�y��������:�����7�OBDD�p'���>��@{���
�߉6*��)��K����l�%M�T*��P��G7�����)�W*��4��Ҳ.8<<���������]��0���K���z���(�TD��D�}��X��j�����/��EDD�f����8?/Z��x���?B,6mre4l�z[[[�`0���{TD*���h�.�k�$"��E�[�����r��0<Y�n��l�T*)����[T��d�9�9��iH&SVDt7T��Q�0���^o���\��*��3 ��ADD?�w""z�z��� 
�h��3\�`]2�M+I��E.�uD'%����9t��dt;�`P�+�ѧq�ݘ�S�U��p��'��E8V���j�,1b�P����r����=*�a��������vZ_(���W_�����ʈ��&S����_�l6ch������ϑL&M���-�>3�]e~~�!�����ۓ��ܻw�n���#qreeŢj���D�95�C4ʋf�v;b�v�'\����󋓆������� ��f��7��� �DDv�D?��+\}ixh�) u��&x�!�f���J4�`0�?�\��y�`u��A.���{Z\\7nؽ�*�kkk⺝���0ub�\n<}����ʹ��ě7����0�d
O�>�á~m|/�>ëW/���2�������k�Z�i<~���K�FC����F�.�{����i9d�L&���s�`0��YJ��n�qvv�\
���,�Ȟ��Z��r��,���Eڋ����-���n�V+ܟh��@@���f��s ^�*��"DD6ŀ;�}|,��{��DFW�����>;u	D'�Pw���l�\66F��p8���L&�����N���k�:
��E���
��)�\.�ץ{����{t�}���'���?~lx����>޽{�CB""����as������=��o�\S���˗/�N�N���G�\������u�\.����C�dyy՚blJ�u��곖D"����/L�X�R�=}"�����h������6��s x���9ք��&�{CDtw9<��������p8�_
� u�e�p'����d�ie�D")�J�I�i�����A�{;����z����\������cQE�C�����T*ZP���2�� @��zo߾�������Agggx������eܻwFާi<4�ln�ׅB!����_}T�RA6�Q�q�=X^^��"{���;XG�Q�ö�d�������R)6e2������5��Z�����
���{���w�7��9�6n�HDd��-��6e��6}��e0���f���svs%D(GaK��t{sss��J�Z͢j�G�4,,����f��ظ�é\stt����*��|>ll�ו�e�_� �a�I�E&��Z>��W_}�v��ě��E<zd|�
�^6�1tq}yy�(��GiwwG츿��(��p�7�,�ƞ...P*��k���-��~���@ ��XD�ժ�.a��|~8���y��Ѿ���_���)�x��]iDD4L|$"�l��y ;�
�O���;!�d7I��ۉ&uz��h�Z妟�~?"� vo7W2����U�9::��D"�5��j���Т��C�����'�!���%޼yſ�	�i=zl8�j����Ev�'""�j����h6��֧R)<y���	���i��z�3���&�>#�75́�5c�B��\\4��J��p`2ibn @(�̞����j�<��;�`���x���`08�����_�O��� ~�!"�P܍#"�,��9��ό����������.Jg%T<�P>����fg��ۻ�.�&��V�4�[�H��=���gmm�����7o^���XR-Ms�ɓgH�f�o6����^��\��\���������q���^��7o^��e�^/��hQU�C�LK$�#Udo���
y2}�|>�v��\#M�����r���F�uß��,)���ɭ�px��
nާFW�w"���>��g G�h������i���`0�A���
��.G�(T�Ms`vV&�f��v;Ud?�XL�Drrr]W_@��0�T*��~d�Ѩ�߇��(��#�i<h�O�>E<n�\�^�W_�K���\^^⫯����sC�c�^��L��C��h`gg[\�H$��d�^����]q�����P�QG�PP�������z�LZ�&�L��$R������h@�X,��^��YT͝�a�
މ�&�DD�e�/���*��s l�1D�H�d���%���G9Q_"����l6�Цۈ��p�=�5���E�ؓ��v�8;���
��auU���a2���£G�Ń�j����}k��O�p8���s��������W���e��ʈ�������o�F��t��D���L�������P#�{�����[P��l6���rM$����Z���P���pbnnޢj�I�s:��$n�J���T	����������R���4��E ��U��;�҈��:����@�>���?�ߵ]n�H�I&p�d�g�.�h�H����nito�^G�R���������V�I���鰃�fg���F?``��%߃�����t�]�}��S&���ĳg/��_�+
�曯��HDDd�^���/�;�G��g������|�VKVt:�x��	4�Ǧ����#�Y[�`�R��eT��=���E�L�h4P���d��N��|^��=�d��hM���Q�1���[2���q3��7 �E?��EDD��7O""k�����=�����.����A nPɌ�Q_8�Ԕ:�Ȁ�9�^/�јr;��kii���u]��ɱu٘�����r������gQE����yC������h4,��>���������߇��f3x��[��
���x�������Bx�!�I��t���[ �r]0�ښ����R� �S�J� R�Y�*���c����ak���������i����#d�h���KB��򹮫?����������DD��U�}�	���h_]Y��i��K`0��ύA]ב�2�K4�Ч�l�V�YT�����+;|�z=d�+���#NF��sh6�Udo��K�x�{�'''�}����66����Ҝ�3�\.^��L�d����1޼y�+""������ၡ��`�N��6��r���#�����"������?�����pZT�}�rYq�A���%�ˢ�UO���ew3T*\\���x��h0�*���L���$��
���� ��LDd܉��kW��W Nqhg��1!��d�vY�P�89���	�s^1���Yuw�|>��4-,,��F�$ҧq��XZZR��v�8<<��"�I�Ç��t���V�޽��&�����p8bh������ u%"""����bww���@ ��?�\�DJ�����J�"���������l6�	{^�Ud_���]�� b�i�*��n�+��R��ݎ4Q��D��V��`45���R�a�}������q3����$"��}����? ����OFX}�$;/�2�J4�p8���)�i�)����4�^��^�K��p80?�>x>??72�aXYY�ө�$?<<@�}iQEt���"�Q�[���oߠ�ᥜq�t����g��boo�䪈��hGG����4�����~Đ���uo߾F��U��������EUч��������
�n6�4���):uq�=}i���vcf&nQ5�"��OM��,��h��m\\�'��	���� ��_(��w"���(�`���@�/��`J@s�т�L&=��&J"����h4P��-��^R)���f��r�dQ5�3;;':�{�5���0??�\sy�;��9�~?����u���|�sN�ϟ?G8l,ܾ��g�C,Y������`d��ǋ�1t;���wSs���0=��ԣ�n_��.�KK�Ud_�ni��M,6�`0hQE�S�VP�Քk���{�t;�j�fS�F��'�����K{�{��q���:���
DD1�ND�� �������@;?xNM����>����!�Y�n��|>?�2�&�������p�\���Q�����,,,*�_\\�P�{���7�i�-���=�z�Ny4|���ѣ��X�j����=������_ �:�������`�ܢ���蓜��bssFB�@/^|�K=5�F+�>C>��=x��9::��z���¢8-�>����[X`w3ɗb�z�Uc/Ҟ}2������V�W�pWeh�}x� �+x'"1�NDt�}��O���!�ؽ]�����h �H^���-�e���DR����:�&�������5GG��:b�P($~�i4H�9�e��W
��}�z=�{��/c��p�ٳ���;;�8::4�*"""���S�yc�X0�g�}�`����|'���)llܳ�"�������@���p`uu͢���j!�S_I���x<Ud?�LZ8��x�e�����B��E�M�Z�ƽM�����s�	 ?��m�
�%��w>"�;��8RP��0�F4逡^��Ѩ[T���R����bQ<Цۓ��w:md��b���uq���F beeE\����z���J�x���ј����[8>>2�*"""�l6�7o^�?�N�ӂ��6��6��މ�fg��s�xNOO�l6�k�ɔx��>���b��9�= ��NG��+����jU�u�����v��ߔ�i��? ��;)	�g ~�~n���� x:º��F�w"�� ԁv�.�q�!T�#E�Lf�%MM�8#�:�ۙ��B$Q�a��<~@z������ZT�}E"�b��5�JE<,���4<�����T*�C�1Ms�ٳg���1�~s�NN�M�����̐�e�����={��!�q����s޿� n�ۂ��:]ױ���\�i��[�Z�����\377ώ�&��0�� ��E�؋�w��"�@j��K{�����Mjl#�~��� ^��w"�1~�$��.��@�? �@���F9��n1iw�v�Rq�eM�H$�ǫ\À�9��E�n�B��j�gaaA�\�{xZduU�޾��mA%����5q�u���۷oxp1�4MÓ'O1=m,ܾ�����S��""""3�rYßϢ�(�={������D��R��x<�w�E�u�\�JE�&�H�A0�tGG�K�n���qMT*�S(S)�� ��{�^�Ba��!�|�Zm�%�=�s�*�@w�,n�Oqx�O"�Ӹ�FDw��@�o��_�� [�ؘt��H$9�K��e�"@<W>��kh4Uc/R��\.�^�����t���lV<��O���F�k��<���-����XZZ����rt�{���^����NOOL��������f���[ �Y,Ó'O��8�:�67߉���q�wGA�� ++��bs�Bͦzs~~Ѣj�G�u1h�J��^c�ZM޿7�/@D��)�3������h	��ﻸx_]YDD��w="�t~ ?A?�~=����ѕF�F�2�#�����DtefF�����,��^���~�r�4ڗnovvN�S���!O+���
+t�YQ
]�i<x$~6-�K�t0�66�avv��ڽ�]�\Y)�I�ݻw0r������G�E�R,Mٹ�\.��u�r	�rI�&O����tq/'��`"i/���"�YT��H��3 "���u�Sv�p8��-^h�p=�`����˝v����D4i|�~��� ~�I �O$�U2��Y�F]	��|�5��8ݎ4��պ@�̎�f���W>�ժ�V�#���MOO#Qwo�fs;��K�B�5�n绮�4�VVV���dh���L�����F!�>��������,�ݻorEt[;;���$�ǃ���*������+++Tbo���ݎr����E��O�ZE�^W���D�v�yu���9�:�JDW���K{�@p�%��[�s���x7��MD4&p'�q��>h���4�4�����@lz��j&O��F�TuDC���l6��48Ms��2��t٣��b1��cv����ʚ򹮳{�(�|>���7 ������*�A��/����>��-����F���;;�B��X^fwu�]�{��^���<b1vH������/=3G8���f�v���}\2����>Tf�f�?�x<!NU���j5q�fffƢj�&�ȂAu����YT	�!������ GX��w"7ګ ��U�}jt��$s8ʀ�L<΍?A6���ѕx\p�:�����L��v+�H�At{R��v���0r���fx�f<x�C�S,�N�YT"�L��}c�W��u�$""��w||���]Ck���ũW4���899�ݿ/���3�7���j~!6'��8���ZT��d2i����D<���"�(����Y ]��k<oH�u]��iUCw�:�����W��������Ѩ]��@��	�/y	n��r���x
�åҦ8�N*�>D32Ηn�������N�]�Rwi]�qxx`Q5����<�Qu��n����wUD���bx��1 �������;�EDDDc�����g� �TO�������ES����1H=�j�BA�fzz�HԢ��Ѩ�\.+�,,,0tg�V���s��?�JYT��H{��H�����h��F��tbjʧ\��4d������;ǔ�H�������@{W�����    IDAT�I�x�w�4~���H[��KT*����˅�i�>K&������W`꺎��S+��D"!�0�d���n1�ǃ��q]?P�{M���x�칡��l6���-�"""�q���k�;��G�#S_~$��/�n�떖��,���32!���wzz�|��N��st{�9M,��뵨�(���t:����V�����F]����{�+\ާGX��Dd����_�����@{dt���H�b���v�n�Q.�F]�Đ^S
�G0� �L)Ç��#��ZX�}h���s�5�B��]�i�a���88ط��r���\.�J���S��w��ԔO�>���זJ%�{� �㉈��jss���NMs������T�^�XDV�d�i>|�.��ժ���]�c��Qvq7S>�G��R�YXX�����r�����Ivq6]�Q,��H�ȸj�:�ƞp�#Y��	>x��m"2�D4lN Oqs|͗ ~����,��4MS~����h!�f3��Ld���Ҥ�8�io�X���E��K2���2�k�d2�@@�9;;�E�%	���iA�����[~�3n�/^�04f�R��իoŋ�DDDt��x�����ϟ���;eA]4���-�����`0���%�*���tq_���22�/���﷨"{�v;����1�ԬE�؋��?==�S�OD@�Q�>�@����z�lI�������L��L��w"�T��g�o��Qu��!pD@6ˎ�DFMO�(_wz�.J%ND���)����0�Lڢj�g~~Q���l�߽��W��{��)�  .���=��^�[P�p8���s�|r(�^���o�F���GDDDv��:^�z���sq���ŋ/�i?d�v����mq���*��|TD��j5�r9�h4�H��3�����{�����,�g ����{�ÁX���DF�z=4�Q�1ּ^���wN _ �%���<�����w ��[""�Dt��x�}z�u�J<α���D�I�)�bI#K�!u&�t:(�9��`�pX���� ;��)O�cK��N�1�4\��kb��F����C�*"#4M���OċS@��7�|�N�cAeDDD4)z�.^���ZM\�����s�IY+�͈�����Zi���� �1,/�XS�M��m�����sp:yy���<�2�TO���u�]���33<o$2�^�?'۝��π;�����_�O|?�>P$"� wˈȈ���\�gFX�!҈�8;�+u:�J�Q�A44M������PP���$�I��|>'v��ۑ��w�]vϷ����y��c��b�`�@�:�޽��Ә�wﾡ�����曯�`�S�����~���qm4�Ç�,�����%N陞�f�5uq����4B��E���ɉ���D*Ő�t]G6�Q�a��������L��S"��\�;�_p�2Dc������`jt��$`���~��@���f��;�4qT�!��#v���|>�/�DE�Q��@]�Q(,������ǀ�9�N�x� �I����b�i�B��3��'��n)���5ONNP��[T���b�bB�������q�v[\�L����nAUdT�u���]qݽ{�t:-���;8؇��}i�]��T���Z�*����YT��d2ꀻ��54��ӟ������͟;�A�z��ς@ �|ΟM�������w"R`����~����qh�9 �d�h�I�}�MA�˱�4�Q��J��С6&�P�[��eH͐L��C���S�������}�{��E� ��͉���2d�D"i(T��:^�~�NSDDDdH��īW��ڳ�����y�"���R+�5^�++��D �F��\N�I9�H P7D�Osz���
����j�*��rM"����vyy�JE}��S=���v�l!�������b�h|x/����ѕFD��tD�t=�~�~��O�wm_a]DC'�׹�$����^��p�F���H���;Y�A��u~~�z�P3��D"Q�t�����n��m($����n�kAEdD0£G����|�b�hrEDDDt�������W��,޿� �ĥ����o�����"�~�E5 �k����/�Ʋ�:u3��9vq7�tv��3e��a�wq�8錀���y����ϧ�|�F~t� ��{FW��D�0�g���p3���=��x�,Tz�
�¨� ��`SS�i��7.�ȼ�c�@ �p8�\sv���f��꺎��Ck�! ����n�rM�X�{��x�x��9�D
 ���C:}fAUDDDt�
yloo��4M�ӧO���,������b�jMs����UD@?W,�������L�����d�k�ɔ��Z48i����"Q����&6>���#�bs_O������[0�Nd��Ms�
��8���+��z�ѿ��azf��j&O�TD��uDA�Q���l6-��>���VK%N�377�|��t���,�ƞ�� ����k��G�Z(
cvvV����akkӢ�H�p8���3x���t���EDDDw���	����u.�Ϟ���岠*2booW���D�L�,�� ���5M��"�Ijn�r��H�ѐ��:���r��wJ�k4�h6�5��Nd�2)�ndB�@?������O ����a���n��U���S\��FX�Hi���R�D��v�`"�qҦ5;��C�đͪ�H��8��>�͠��ZT�=I��vo���i�ulT��=8���/<��G�#�;��ln���""""��vv�Ŏ� ������Sh���%Y���bggG\��q�,T�TP.��kfg����Z�v��:�Uus���9�����{?����a���K�p����n��R_ ��@ �|����}���}��w �����/�l,���1�dJ�f��W��'#��h�8극�8��K��Q"��z�՛LҦ7.���+��9��xI���̢j������e�\^��Eó��(�4�MC;�kk놺��j5�~������hh67ߢR9��bӸw���l�rI����`u�}��txx�|�p8���hQ5�$�E"Q����t;����A$�����لBax<��!�l���v��v�_Op'�!����� �`��h��h2$����7`ډ��#eyC���V_���l���hpR(���?w�H����*j��E�����
�\GG�C~��c��>����^���H�H$��;R����˗ߢ��D
"""�^���/�E�)O���_����U�[[��u�g����Z�T*��?����j�l6#~g�����{i4bs�DB=�w~^���rM,6mQ5D��Vc�]�=1�N��D��D�)��q��F?��K��`�	�� ����;��T��9�Ƞ�i�fu�P��{��Ba��)�ѨrM:���f���B2�R�)�Vy��*kk�p�\�5�l����#Y#
�ѣ��^��W��E�uaAUDDDd7�v�^�Hw��}D�1�"I���ёz*��i�o1��������������p��s��]��g�H$~:Ţz�_:3 �>�e��B4T�� ����;?4�~�$q��g �'�J�IT�1].�a�eTɱ{;�!������f7.
���)�0�n�~���<��z�f3�dC��K���t�O��Nt�n���UD*n�O�>3�x��-*N!"""���u�~�Rlԡi�<y���)�*#���\\�/AF�1�� j�|>/v�^XX��鴨"�9;;U>w��l:d�lV���x��<l؊Ţ����4/py�B��ucM
�sb(�'I �)�߀�W`^�h,0�N4�c��hȤ����7��<�DFD"e�^]�Q*�-�����Mv�6��ib�7�ˢ��XT���\.���)ה�e���[Tml�?W���q2�x�z��ڃ�}^�!"""K�E�����n7�>}���Q�������ml�c�jI�].7R)���^�R�����[T��4��g/���J�����F(��"���h�/�ٝ��W�?��ϜDÓ�3 �G?�wމF��pD��f���o�
��o�hȤ�;��p'2&S�=?/��e�w����Թ�ngff�:*u�O3?/w�c�v�$	D�Q�z����c�*"���{������7� """���.���C*"I>���NM����hQE��e�l6�k��L�y��3����'Q�D�d�H$��i�:��U�Է�i�E!Ma�;���W����x"Ӥp3�~�~��? <a]D��P-�9�
��@���iܕZ�;$mRK��4�P(�ϧ\#���H���;��H�XXXP��ժ(���c�Á��{���meG/�F2�2.��jx�� �Έ���Z[[�(�K�T���2��Ζ�Yee�Ǣ��M�u)��|>6�1Q&�A��S��Ľ%�i/��v#�/|�`���9����)�Q�@D}�����%n��FXѝŐ-�p���� ��@���GV�MI��Vc�v"c<���rM�X���H$��ۛͦ8����x�R�.�4�TR�t�>̧�Y\\;�
rWG2_0�Ç��u���x��t�]�""""�I�u�~�
�ڍ�{*��F������Ӊ�U���N��n��k���,��~:��x�0;;�.�&0�*���=�p8��1"I��.H��P>g�����U�}7﫣+���`���v���@�o���َ�h�T_�����/�v���G]�D�¾�V��M�H$��ٽ��TJy ��=��i+����!|����x<,//+��z;;;UD�r����38�-0]����+�Z-�*#"""��v��W��E���p�i�<y
�W}�̷��'����
�,���z��x� �"[T������x�^D�1���iO(�H�r��U�U�ۗ�����:����kR��������n�WFX��b������ߑ��v�1'�Wff�U2�
��Nd���zs�]{�/
���Y|͐J������p�C�"�'F�S�E��7�t��k����l6,��~X?�%�o ���6��5��j5ln��y<<y�a��t:88�Vi�ظoE9���DyI�����R����v�=Q�ۍH$bQ5v��X,)WHgD�W�s*���Ԕ�����H\����g���RBd �݈~���h�;�ߡhg[�1&�LϨ;.۝����ib1u��R�`Q5�!]Rj4�5A D �W�{�����n鴺KG(���KXT}����^ �L''�TDDDDdL&����.�`}}Â�H���D���D�',�����Kd��D"a�",ݎ�?�'�t:-��>..��V��5l 5|Ţ��?��ш$����i|>������:���x?D?��G � �8º���D}ګ ��U���\Dw��J�R�Ng�e��p8����纮�TRwo�����C�<'P��H��T��(�q����)߿-����`roo����FcX^�'~�JDDDd���Cf��1]ױ��%���؀��h�
�MӰ����Y2��r�����vr9uw�__O�����n�8���p7��W܉h"�����O �px� ~`&�d_�+`����Pm�bv���G]�D�^K*�s��ljjJ�"΀�4$��{&�������u]��1�O[affѨ�#x�Vc7��x<x���ص��n�իo���,������8]����K\\\�k>|��)�U�ǔJ%
�.�SS>���YT����uqJ���<\.�E�K�������N*5kQ5�"��_����m�s��4�%�$�N���Q�1����9�h������ ��f���<ɖp'�p�*��W ��s���4MP	��z�V4y
��-�q�!N�0�j���\,�;3��E�؏��A2�T���h���}*������m&���G�����(W�c�ƈ���F��<�˅�O�����(��l�����58�N�*�7�������,/�%��(��o��5�M4�v�>�,@:K �>vqW���w6� �����x�:��t�]�>��+�_��
 <�҈�LR�Fn"����H�v�
�;���]4����K��:fH�����:j��E����¢R��i8R��8R:�ϡT*YT����5�b�.� ����r��+"""�Z��[�`0���{TD�l6qzz�\�v����dQE�V*Q���+�3��\.�^��X!O�ۑ�H�=V�p��p��UC4�pW�x<��^x%��>���
W�w�`�h��
'���yk�K �G�E<2�҈�J�ft�c ���&7��_�������%�C�r���?��9�b�N��9?�f�v�8q|}�\��8���)�躎��]�*��Ű��,�+
8::��""""��8;;549k~~���;8�G��V�YZZ'�p�/�{�S�����{u�ԬE�؋�s�B�?d�j���_�5MC,��"���3j���W>��="[q x����/���$?|Н��;M*n�s ^��V_���Ͱ���3-\��:���fff�s�N�r��!���ud���t{�Dn�:�����XXX��;�\svv*�'�x�^<~�T<Ĺ���۷o,�����hx��6}�|��|>���t:8<T_�t:�XYY�� ��f3h�Z�5Uc?��z�( POJ��U*\^^*��b�p�.N��i"��E�^o�e�5�_p'"[s��/q�9���;��Db��&ɇc6��9f�� @�����B��\"#4�bR��`Q-���]��"t���&u�*���A1ݞt��h4P(���l.������n��D?@�Ç��v��}뺎7o^�5�����Q�����/��v��N�w�x8*''��w幹y^D����8==Q��Fc��Ud/�RQZ�R�:1|��_$���3܉d����d)��E���X��w �@xt���-g��y ;�
��SeDdK��)��C!�~�ѕD��!e�N�u�J�n-4��!^*(rUc�Ѩ�bX&����	����{K''� �am����\�����xhO�YZZB��E֝�mT*�TDDDDd�z����w�P(���U���������\�i���-�����N��8��n]�'��R��$.��W���r�,���R������.a��|�;;��������'�����7�i,1�N��}��� �q3��+�D$�6A��p$�;�����V+�;d�XN���u]�
H��^y^�2����p��튣���y�^1��n�qttdQE��`0���5q]����R�d�f3H���u����e2O&�Z�D�0�ě��n#��*פR���Dj�`���T*)'~h���i�����%j��r����Dv�h������?�8��!��P������J#��w5���#\����h`b���uJ��9;��D��������y�\B�ӱ���FD��9��M�v��H$�k��3t����muu��/� ���>#�t:���h�z{���o߾��*""""�mmm�!:@ãG��S��<��cooW\g�&}��c�eW�ӉTj֢j�V���=���^�'64��\ip�bA���9�d�;�K�.BD��a���
�{GW��d�u �@?�~������ED6c�]�PPo�Q��A$��U*�,��.4�̨������qd.���gnn^�rvvjQ5�����C����.F�޽����:�����W��BDDDwJ��Û7���y��D���ZT}�Pȣ\V�E�1-P�UQ�V�kxTi��{<WNo�ۑ�Lgf���4�5?��)�����xi?��hH| ~�i�����4�g������	���ˣ+���*]ו�c1�U�����2t��v��2L8���Q�)p�dRݽ���R�E��i���kJ�����>���x踷��^�gQEt]<���윸noo���DDDt'5��l�������Md��]vq'''��>�/6�    IDAT�/�!��(�o�N'���C�P~�.D��i�4���s�>���D(��"���h4F]�X�:�K�	"�[�������-��w��>�-1�N�t=о��_�����."�	զQ0�v��D2iÿ\.s�hȤíj��V�eQ5��H$�ϥ�I����8����kNOգ����|~��V�!��YT]��z��܉�\.���Ȃ�����F�������tcC�|C�V+��(�`��GM��e�n_*��ϳ��Z���r�����q~~�\Ë����P����A$c�]M�\φ,Dd?�����f��� ~�=���.a��>���;�hg�	"����2 L�{�R��G'���̿�ᛙQ��{���!�|>�l6cQ5�3?��|�j]�R��֌uox�c<x�K�7��t���[�wDDDDwݻwo�j](�8�N<~�D��K����/����X�l�^ggg�5333�s��L&�|�M��rYT�}H{���+N����;���K�<���)e'��L@?��; �4$|G�A� �� �;�m ��
����.""�p�p�J�os	�N'�a��P܇���(�y܇-�Tw̺�h�Z�ZT����~q���)��, �H(�T*�(�UD���/�l���Nz��No޼�'�!,--[T]�h4��f�kB�0fff,�Ⱦ��Ԛ�ann��#��)� ��&�&Hx�^�B�=o�tF�D<%���LjRċ�D4��x� �����E���IŇ��/�� �� 6FX��b���N�D�H$M����N��Z�]%�I:ؽ��@�^�������^�P�nO��n��}�~�D�{��5��SSSX_��#NOO��񵊈���������#q�����#rp��.�c��T���y�OM��vŋ≄�������4/�S�RA����s�Áp8laED�����j������C����� ���� ~ 2ºh���9}h��� (�jT��N���FH:�
�P�H�d�����QvU&�r�4b�
�������p ��U���h�/-�Ȟ���x�����;FBãG��t:���vvv,�����h|���R�(�hZ�3û�k6��d��5F��Ч;==Q>w�݈��I�Ҟ���4\.�E�؇4���K�u����k��"6�R��s
,M�5 ��/�ww� ~�#���` L���8�� �/ ��,��h�і>�^/_�T���N$2p�aq8�F��5�_"�>Ho6����5��D.�K�F:��Og�c�����Ї���t��7o^���x�4"""��J�u�}�F�,�����jMQt���>t���؀��R�iJ�"��r��,3f(�ʳM�x��Ţ��'
�b��IgҾ7A|��;��;�D4a��gU�~v���S�,�������ߡ=�O ~
@�� "CRǡ��+u:T���NDv�r��kJ%v��h4�|}�v�8??��"{�FAg��*���9��y�Z�1ҧ	�B��Q��.����4~�kk����}^�!"""[k6�ݕ/d.--#[P]wqq�tZ��=�����I�c�(����hp�nW[����U�U���>�4��hC&M����:"�c�]���*_Gt]��&"�T ?�U���C?�kН�w3�y�w� �� � �=�D�4uG�(7�J�oq	�Ѩ�ݾ��!�F��ee�'\8��ԔrM.���{����D"�5gg��n6c���,����4�=dj�*��-�����h|���X,*�h�����X4|��~���*���\�LZ�v�avvֲz�$��*��b�p��M|�t]��H{�4�Z��N���������l��Z ��H
"�	�𿢟q=�G ?eAd=�\ك������������!��V:�Q���
���������'uoo4����R��n�+ ӧ	���N�P`�XZZF(��.������kz}gk��ݏ� �Srh�Z���N�k�� ��E�S��A.�W����c0��B���/h�����6i/U����.N �������j�������G]��B ��?|�����"��w[�o� ���ڹCDw�d�hE5��ɛ��f5fjj
>�zt��׮a���#�s9�͠i�R)�l6�<��O���*�98�7�����ceeU\���˱�DDDD�\\\`{{[\����p�d�vxx t�����i�i�E��ˮ�&���b�:�T7a��I{���`Тj�\V7�as."��Ԥs4"�;����� yD3M,��U��x ���NDw�*��r��,�f�%Rr�=ԗ��j��1��l��lZT�=��q�%����p�=�5ҡ;}�ߏDB�.�ϣZe�vkix����U�r���c�j""""�������JÃإ�b���8=U��O�b��L�rY�_�����{��ԯM�hL�+��\^^�VSOf����3LҙA0��岨���l2�"�{��E��L�/l�+��y��p�[^ �3�-��x9����<MӔ�h4��n��j�a-"��J��b�zȤ�;'O_"����h4P��-��^��ԇ��z�W�jyyҰ���}Kj�+���D��D{�.޾}#Nt""""����M��m�@ ���e�*������Q��
�)�>S>�����a�z�
��rR��i����ipR�|iO�S��qyy��皦!aw"vpW��R�u]gN������g���$��z�ת����җ���L��s3GB �2*7&1#�M8���IB��$dK� ᦨ�p�}�!��ٲ�N ���L_�����~Y��с����Y�Vu���yx�a��ך�յ~���}_�� <���Cvb��dx�|�� xԗ�<CJtL�3U�7�Ke6	2�s�\fz��t]H�14<�������g��2��G)
�P�V�S*�����PE �P��)���O��B�������x߁g ef��:���\�J��C�tzVV���㚦azz�����0���^>_p��BCR��mV�T�ץup"�k6��V�u�PHy܉ȃ��+ ��� %\��c��޶ ��� ��A=KZh�R�)�Di�Y5J�I����|���@���`E�/�L!
+�a��hl�:�~�3�����A�"���������Q�. ���
��N9T�޵���b���G�u�{�y�6��N�8!6m1�}�:�66ԍֳ�sU�-kk굦t:�@ �P5�P�n���Y^�4��Q6����"�3�v��2�Z$�>��w"��el��3�}c��ޔp;���	�zח���2\�S�;��.
��Clp���Ԕ�z�R�aX�0��I#���:���C�x��i�4�[+���u��{����w��Y��:m��U(L#�U?���O<�PEDDDD{�w������>�<7�F^'��-���5OMe�H$�țVVԓ�"�S�G�T�@��n���i8�i��H��Y��w��y��H�l6�.a�E"�K "w�a;�� W�\����(�[<�] �1�DD �Mq�Y��w"�TJ�i6�L����TVy]_LÓ6��>SSS����e�&;�������e��;+ଳ��;~�i4��""""T���SO�;t���B��~�P����3�}�J����'����!��K�4�rY��Kk�4�f��V���Gڃ �:��I�Ҵ ""y����\�r-46��/� �s�"��a��X<���`5{K��C���vDc-�L*�3��^�PѨ:1��'��D�ϼX\w�o�6Ǜ�&*&�������>�=�Z���:t&���z����UDDDD49�����D>�g�y�C�ݴ��^Tޓ���qkpTL���ʲ�|>��{v�֜2�)�|dn'i�c{}��;I�{S��C��MLpW��P�z)��<�% ��� 
.�B`���;�C��p����)q3���J��S�D)=EZ���H	A�V���6�����V�zݡj����?�Lo�}�����Ǐ?�L1`{CW:�a�&��;,Ѯ�x����&�|>�l�	�N:q�i���/8Q�gm7�[�g��<���V*���$]ב�d�h��mq�ojjʡj�A�CH&��N��w�@  �I=DD���� �@��D��o���^ ��awK!"O��)���lpW)��<M�����t��MNA����[*�G���Q�Lo�B��\T6M��+V�-�����FŢ:E��i�:��'����@EDDDD���lt���3�f#����G��<����>*�V岺	uzzơj�����٬:���'=o��n/i!�H@�9��Ȋah�[n�1�����SAD�ai ����ܱ�թ�� ��=�	"�]c��Z��w"�d2�\��t�h���fMӐɨ���]N D"�T޳���Q���V^/�6��t��{��g�Ɛ'�C��G�ڷo?���V��T}"""",.�@�VS��D��p��� �?���i:����P5�$4O���BU���S6�ec�ͤ5�T*�CN6j4�v���5MC"�p�"����l�]�X�D��DD$:�C >�����L�K�� �@=����`�ꦣT�c�T*Lp'RJ������+�H���h��L� ����9�H$"�^]]u�oڿ_��j���ƿ��!�q�A�'��_���TDDDD4�L��w��8����l�qP����Mu����|>���J��.�sh(��ix���ϣ@  ���p677�?뺮�k�4�jU���ϛH��j�p����&�k �� ��/�c���� ��Z�!"�+T���^f�&*��	��I'l��W:�No�6^hx�\Ny}ccC<LFÓF��z=&�P6�E4S�s��"�t�Yg�M:kk���z""""\�Z����]�q���8T������)i���>��u�=33�����tP�V��HkX4�4���t:�P5� �%�����a��T�0���h"D�� <��Zlp� ��A |;'"��i�ƣT*ű�
��z���e�-MӐL��H�+4iӄ����u2�g^,��z
�������Gh��y��^���u��'�� �W�����8v�I�*""""�cǞD��Uޓ�L!��;Tml�h4����/p�{���j�h�x¡j�CZ��������*���pKp糝�J���~�u��%���� ����A�k�4��x��| ��Inp��J���v"�x<�L������jV4�4MG*�>P������@׭��@�\r�"oH�R�D��{��tڽX,.�Y^^��h�`��O?������|>���3i�����d2��L���m���'�u>]G, �B��o��h�Z �z��~��0P��ھ�i�R��\.�R��T.�R�l��\A�RF�\��$"�^��cǞĹ瞧���3�F�T�3�!'O.�sε�����Ĥqڝr��v��P(dy���4j�-��|E:t���p8�X,�z��`U�MjpO$�������d���-�]�9���#��g��B��E�׃����躎`0�N�����:DDC x���_ ����x��#� ��v!DD{��R�w�2��������j��6J���f�~���-��bN6�N�bC�hH��[�67y�cT��M�ĩS'�����/�����;!"[��~��΢P( ��c��<���1����o�>�f7U�U,..bqq'������X[[œOC��1�DtzVV�1==�L��B��_��O?�`e޵���3�8�`�: n��y6������U��[�?NOO�ر'�6h�F��F��h��1�˳��F�Z�n�@`�뚦!�Nacc���&�a���z&�}g�d�?�D
�V�ST�ሲ�����N�s<
�} n�Mt���y�x �YnBD4�R��T)���HE���#Ei8R�r�Rᦡ�4MC6�U޳��M��4]�����P5�
��ϫ?���U&�;$ba�x������D4�`0���:�s�9��{�8t�
��c��.I&�8���q���?�aX[[�Sǎ����O<�'�x�����������=�K/�L��2?�����L���1��K8p��{R���$�U����ꊲ�="��B���_;ml�Z��lǏ?�\AP�T�k%�t��6�V7���T
��KVD��4�lpW	��ܻ$"-?�� x)��8�n9��w�h ��� �c��h R�K:�nN��2܉����M.�Inp�3�N�d�2�i��������`M��o�~h������E�����#�WV�Q�p�Y�������s���9�\�q����'M]�133���\~�?����>�?������x�����X[[s�Z"gߟ�����=���С3�?��w�̻N�:����������1"�z�z�X����i6�۬X,*$	�B!�Q�R��>������U+��y]��p���G�.���+~��x+�O�\�'���s�Nm�ۅM
U�{ @4s�����ns�H!#
Y^7M[[LȲ����H�S7��h/)��Z�R����)f�׫�*�~�χ��9�=�J�Z͡��-�cfF�����ر'�������y\r饸�Kp�%��Йgr��|>:�C���~��~𿯯���ÿ��c��w����G��s�R"'O?�
��A���|��T�$�;���`mm33����ry��a�����*�np�������]j�j��N��`�:'.��ai锃UM6)T$�!���:T�d������� �e�,4�M�Kk�HXy�0�*!"�$�?�
 o�f�b���=�� X�B�P4MS6��Ri��{��L�&����un^�(�N)�z�.�Nm���י�n?�?�lvJy���C�xO�0-��/.2��)g�y�ؐ���Os���B�.��"\r饸袋q����"I-������8|�0 �V�����6�������c�����&I"���8v��;�9���:�<�ؿ POפӷ�x♃�;w�4��sx�)NE���U<x���E�ud�9�������fg��Գ�,�m�h4�n�a/R�4��uG�T�n�F�h��T*��u~�D;i�Z0M��-��e������v� .p�q������z�{ ����P�w��Sa2�����Vh8Ҩ��g��
���( �i5�|�f}��4���9X���۷Oy��h�T*9T�������è�F�D5??��/��_q����#�d�Q�����+q�W؞����=�G��Q�㣏�;������VWW07��d���O�YYYv�2o��{�Ԕ����9?�49G��i�R)#��>�^(��n���ue�{:�������Q�R������t��v�V7�k��$܉����V��H$�v)cI�4�!�����;��h$x�� ��r-���	l�� ""�I'��lpW��d�;��4����%5:�P��T� �j5�h4��;������F�i�#�J��Y����'��4���::S���'��D!"��ø��Kp�3M����%yZ(��Wl�]���ɓx��o�}�<��*yēO~_|��C��X\�t;�<��|����d=*�����L&���6*��0�>tݷ�u]בN�yH�F�JY���ɨ�Ih8������>�� /"�f��w�H$�lpg�=�Ȅ ܅�4�_��v���~� �"��.��ȫT)ClV؜Kd�����<$b�ߏx<���R);T�7H�� �_ '���:T���۷_y�����w�������{66�|M�T*������/=��.�L|.�{��ߏ#G���#נ�n�_�������_��M�j����U
�͎�@��x�cV�M�r�z]9�d���lp�bq�q.t}�l��#��s����@�RQ�_e2S|o�Q��^{�FcC�t�U4٤��x<�χ~��PED{K�� `}����� ����Z ��K �hb��/��`sE��    IDAT;�HI���$T6�lp'��J%�	�v�6��J���w��A�^w��ɦi2ub>7���?��G���`E�������,s���@ ���{L���O>�PED�D2�W��U��c��[���{���糹}	�Bx��ĭ�ކG��(������ѣ��bc�$:v�I�;�����BU�m��K���x�_F�ߗ�����C�x��6%�7�p��Z���i'��l���X^�4��:���Z-�tr�~�;��" ��Un2)��n�7�2 �"����}��e/��j�u�n�A4��2��< b'is�\f҄�R�4|>�!^�i01
���z�����������=����"d������CO�<�L
M�p8���~��n<�ȷp��w��/��@����4�|>\r�%����������#װ�h���m,.�Pޣ�:�8�Cy���ܞ�}��9T�����)�g2S�~c�����h4�>�Ik��dBNU�b��5�@��IA�a8T	��%|�Mn2	��~�| >���wk���i��lpO&���^'�?$�dR}V����ɨ7G�lm/)a�R�d���� R)�Ai��vG�4���)�)�6�P�p8��9u�M��������FE�u\q��p�]w�����G��F0t�4��7��r�x�[���}W^y%t��D{���	1!szz�X̡�����cuuUyO>_@ �߷����>��i�Y��0N��D��n`�{Ik��DH��#�QyY���yY(R�I�z,���v:��� �2=\i>=	 	�z�!"�
�y=���f�͹D*�:u�Z�:T���F8��%m�Ic�ix�|A��e�q�;�\�PHy���)������O?�4z=nN�U�|o��:���_ß|�8|������?�R|�������nx'���0�0��Sǔ�h���9T���:uRy]�u���:T��l���������m4<i������`�መ
L���	�s�H�0�L�41d�҉��: ���]�o���� ��ۅy������>�
ӧ�,E"�Ha�0P���h���i ���v�-�5���� b���rY�aKÓ6�76�:"RC]�������q
��f��KUDDv�u�_q���43��ϻ]����i���������Ç��s�)�^������-�=�l�z:��F�!6����q��H��2��rM��'�Q��6�٨���PO��&��j�-e�r0�a"��I��}���W �G �q����o~�s�� \�v!DD���lpWڬ�GyY"�No��j�g#�y��v{MMe����6���C�xC0D*��9_[So����b1q�ui���8t�L�3��c��wA��d�9\���Ϳ�{6.��B|���o�;����.���p�ؓ�=�1��	�N�'P�Ba�ݟvgcc�~��i���V4���2���k.4i-���}��t���^��1�]-��"�1u�� ���B�6��j � ��Bj~I�8�ϊa��R�>$�2i�'���K��T8q�N�&�4������i(�~���#233��nVV��ƻ��42�����*��u�*"�ӱ�p 7�|3���o��_����K�=�P(��o~�������8���.��P�����D"�|�ͽ���Q�fg��B�;���M�o�^�a`S�F+�o�p��X6��K�k��*����b�����NDD�� x�\�cOa��p^� �FAD�U����Ǚj`ek��L=!�:)E�M��~^Ǖ�lnr�]4MC&�N�.��hm�|^}&�X,���h���iu����*�ݮCy�vz�ړOʉ�D�K/�w�u7���C��ڣ�(����W�_���Ɵ?�\}��8"�h�m���CG�8��-��i�X^^R�35�E(r�"oY_W�M�3�U��Z'�KZ��Fc��U3���&�Yk6��"%�s�&�� >	�]n�W��}po �y ��!"r��+�C�����f�͢D�4���L&�i���n��f��`E�-�L*7�L���pB�R�T���5���|>�@@�Ẵ�n
�ӗ��Ĵ������GD��uW_�"|�s�ç��>|>���h]r�%����K_�9r�A6��Z���5��K4E�0�PE޵��Ӵ>(�i�x��vgcc�~��i��rV4����X,&6���:��8%BZ��1��h���>�K�`����� �~濓� �.l���]��I���$G$�lV��Nd%�*�v��>�B�Ez^3��^R����&z��C�xC.��j=���T⡂Q���S^��k<��*������:�P5D4(�ߏ�9��������/r�$���;��z+~�kx��^'V#"�=��1����3��>b�NŢ��wvv���a�ņk6�۫�h��R��NMM9T�7T�=$��٧^�+���~D"+"�[��^����wj~g'"o�`O���4 wa����Lz�J&�h�Re�(�%i����P��K*���6Sh8��z��\V�|��e��M�bq]��G���ɤ��0�}���<�������u�*""���8|�0��o��[o�ss��BD�23;����<����ȑk89�h��Z-,-�R��D��;� �E�;�$�t:��]6+��kVlp��:"����L�D�����)�D֤�^'M8a�;�X9
�K x��ܭi >�nBDD��T���D֤�b���I$1��>~�_l4��h8~��zïX\w�o��
���ڪsy���P�a�&�ڑj�H����n8p�품 l�N���[��׾�Fw�1r��q��}�=�)��z�R�,6u���:T��ll�`��t]���p�P�t:�&=Ik��D��xm��X�'��f�	�*�pHy��;�����| O8�o ;� ��nBDD�K0�ݒi��b����Nv�Ţ����#�!������r����V�9X�䛚�*7���>�岃y��i��Q�E������9T�7
�b�C5��KLY"r��i����_�"��n<x�품v�o�>�r��˯�^��W�ѝ�e�n�N�T��1;����2�����#��#�^{��1�}>�SOt���e��A�hp�z]�n��:	~�v�ܹ�Id�k�jR�;���; ��;lp6�G ���B���G������k���z!���4M���n�TJ=&{k��畍�i�;p��Fk�I�٥R�?�#��f��i����ƛ4MNo7'Nw� "��O^v>��/��ދ�����v9D9��3q��w�_�"~�~��r�<mq�xh����un?����r�\�t
�V��bQy}��;SQ����Q���e��/�)~�ɤzj!N�sH$�|�Yh����ܥ�""rͥ �`��B�	W�~�� ��v!DD�l�f�`0�PH���e�M6�Y���ʍ�^��4I� �(\ܝ�i:���k�U�-33s���f�������iD�Q�=��Kh��UDD?lffw��~�������w��]9�9���~�~����aaa��r�<���)��`�����tz��$ο����(*���~��@éT����4?o;U���T��vi4Bb�O\g!�~��n��vcKJpg�;�Xc���a���O�I ��v!DD�lRJA"��viQ������z��JÑ6A���O D,S�#m�p2�4|>��u�4Q*������x����i�P�c}��� ����߆�}�kx�+_�@�/|�����>��n��z����E1�}aa�)�#������Ő䚹�ݮ�p-Mv��H��T��qm$��� ��j5��'WYc0��`0��.�w"��w	���\]ڦ� op�""� 6�s�GiSXt'�2i�OJ�C�h�MN����`�n��l6���Y�&��f��2#0==���h�VVV��{��"���S�N���8Ti��Ç�}o��zN<�����q�G�G����s�$"���z8yrQyO0���CyS���nW������QT^��h8��U��}��>���9lT�Va��Ӕ����O��ڒ���<D^�n��]%T��0*�ػ�7 d�.�m����`s;�X�ܹȣRR7��Lz~H��48)��Ѩ��c�]2���z���v�I��Ţz�vgzzZy}��:=����>�MPDd����B|����λ�������T&���7݌�~�A\x�En�C�'O.��w8�T�2M����{
���F�X\W^�Ü0b#�4ĉ��z�g}�j5�=�/N
�a��5&��IA��ND�'\�a ���U�6 ��vDDtz���j����hLy��#m~H#pi8R��4♆�H$�Ec)卆����VV��ƛr�b1���S�N����n��x�����}���9�.�g>�Y�r���%":}�~_Lq��(ԇQ��,//)���LMq��ݚ�&�����۫RQ�4Hk`4i�6���mi�!���&��q��ĸ�C <����o�o��]�>�Xk4b��W��qeJA��A��v��ɖL���)�`�HTy��9H���ԛ׵Z��2#0==����vP.��ƛ����Cn~"�����?�կ��]���v9D��4G�\��>��x������M�S�N���)�ٞ��t�Qi4bsd��~g�ݑRܥ5�ҐL��l#)1�	��i�Z�@ M��`"��Z�Z(v�""��� ���������� �r�""�i���Lp�&-Fy�������|>q<3�W��dԣ���&Nl&��1�}4��������HڽL&#^ZZZ�aK�J&����[q��?���9��!�B��=�󮻑�f�.�hb��}�:uRyO4E>�F�QZ]]Q^��U��;~<�@8��2�lmm)��ΦkI!$�h��I���I��n��~��vcKJp�9ў�3  �t�6��"�O��DD{�a�ע�(�~����-[U6�Y��Ջ�U���M"���ͦ�M6i4��|E�	�È�ԓ�E6��mj*#.�K�tz�P^7���D#t��a<���ȑk�.�h,>|=��8r����ɓ'��"�;#���5��^Mӑ������-t:֩� 05�CVv1M���I��:���t�j��i9U�>R��C�e�6'0[a�;�Dz5�{�.�i^lp�Y ��NH"�=Bڄ�B���8F�eRCj�Vs���'&`z���M�r��v�6���j5�>�����z�Q�s|��ɔx�fuu�MD#P(���}w�u7����.�h�%��r��O|33��D4�^����S�{��8}G���T*)�ޝh7L1ŝ���U�H���S��:��������b16�Yi�8��J ��[����Ƀ�DD{ӯx��E8�k��x@��B��hp��U<������v�i��L�#1-�>�HD�-�^�p�M덍�*��χl6��ge�������n�&O8T�w��%/�_��Wp�UW�]
ў��]����_�e/{�ۥM��'��7`~^�ݑN�4�*�J!�8T�wH��t��ё�&I�|̷�˖���w����=��=6���f��J(�n�c�;ўu��p��x�z�C RnBDD��c\HSa�;�΢Ѩr�����a�]�w>��#%V��uq�6N�u11���������h kk����5�H٬:�smmͦz�9.㦛o�=�|�����,�H�?��q���F�.�hbt:��,+�I����wڽ��"z���Baڡj��\.+w�|>$�ܖ�K�VC�۵��i�i~�v���L�K��R>�}>"u�	�W1�]-R?;��ND��}���.�	^ipO � �nBDD�c��5��Q��]�X�F{J�)48�? &��jlp�K*�np��h8�TZ�hm�8F��7=�nΨT*h�yHiT����xܙb�<��.������ڣn�B4^��W�+�׸�K�.�hb�8q��Nq߷�[t�b��u�=��3U��a��o4iMK
 ���j5��iy="
9X�d��"�q��	�j|NM4��\�v!��w?�����B��h4�T`/��R/By��hOk���"��m6b���Β6�+�
��P5��M땕���@ ��usL�XD��,�N��i8z�(��gq��A��!�(������i\�ۄ�0D4�v����5�=�|�0hGeuU��D��<�RIy}jJ=���#01�>�a���|��Gڋ��z����ns\��DD/�+ �r��Q�B��� ���"��h��S�I�ˤ1�D^&��0��>R�������Ć���M���i��\Vov�����r|�a���Bڽ��}�uu#�ɓ'��hrMOO�S�ߏo��@��r�&����[��������[D$[\T�4���w��T*h��)��|ޡj�Cjp��b�x��.RhC"��{��������K�����hg�i���]�ؒ�y8��h"���>��&��& ov�"":=�a=�6
!:X�޲Ue�(�iQ�Vc�]�46��'�R'U5u.��(
!�*�)�6��;����z�XD����Q�uss���lmUy���4]z������.���.��.��R|���˯���R���z�.𝝝���w�"�Y[[U^�ޥhx�F]<X055�}�k4�u-Mә*n#�����]��)�����m��a/�ٱ���hb<�_ �������J ��]�U:'�E�V�	�D;	���4�h���.r�;�Uv���tj�l6���j��h4������s����P5�3==#.]\\t���t��5��O�τU"�e2|�����N\�""k�wA�χ��9����](#�dC�ݤ���z��ZU�mIk48)��	���Np�n4��< Fd��n�]������I�lp'"�(W���E�¤6���S������<Cnp��
܉v&��7��\0�j�\2�w'e2S��Lo�_>_P~?����xڽ���+��Z-��UC4YB�~�� ��z+�\���p��ć����v�\.=Ӥgm߾�<H2"�ZM<d�w�I�SS���HZ�b��}��:�zB���G$q�������l�S�c��C��-lpW��a%�ζ:"�	� ��vv���T �o�DD�	��D;���HP�4��Ѩ�߷�(���|>�g[J���i��LF=f��������uP���)D���ԓ'��C���翀_��W�]
x�_��=�y�y�Yn�B�'-.�P^�B��8�dT�w6�ۯ\.)߃|>�H@��ֶ�?k(�� �$��/N����"�b��Z0h@ȽDD��| �K�.�N����4 �<yܭu�]�Z��"���N��1��|(����%I�bd��A��t��ɖJ����{�T�V4�����Ķ����Q��S���z=��,;T���/����s�9n�BD?�����������D�9bmmUl4ڷo�C�x���
��lm�~�/��OM�'��බ����~?b���M6i�So�#��p?�hg�6��U�Au�;M� r��LZ�� ~��"���9�8Ϭ�i�Ț�,�������������6�+�MN'��vҠ�!�^��r�����ş���%����ѣ��ޏ!�d�!�8��b���q��os��=�4M,-�RޓJ���;"�z��:�A��E�+�6����n�0��DⰏ4%�	���ܙ�N��N�É�
R�;M�) _0''���5 np�""���BOpA�J��D;�4Ѩ���?v��՛$48i�NJ��d2��iis��W(��76��7ڽ��}�	�i�ԩ�VD���|>��ݿ�o��>I˳D�G�4�������}��~��!�3������sssU�=�d+��0O:l���f�I!RNNp�+�hpR���TZ~�D?�4Mt:��[�܉�<�B ��]�&e�' |
�FOD4qT�>��p��j��Z���D;�F��F�n�+�Ҧ��ô��N    IDATa֋g�i�^W��Ѡ41��	��	���e�$n�P($�X[[s�o�u33��{��"w(�➏|���׻]
�կ�%�w����D����bmmUy���4�~6����هB!�RL]�S�VC��z'ҐN��g�I!lp�O��@�׳���>D��V��~�����|�D�VD�wp]Қ����{"���z ��v�k�� >�	��'"��z���bL�P����J���v�H#jk�Ӗm�Ŕ������m��Mi�� �N��7l����{���C�xK�0-&.-1��h�|��٧��^�v)D��_q����`v���D��&��333U�-�FC|'�ޱhx�rEy=�b��]��p8"6���0%i�W�����8�Z��n�]��
�	�ܣ#"�x�J��8����Q �q�""��4�=S'�z܉v���c)�PqK������*L��vI�3��l��_.�S^/��3>"ss����:*u#g�}6>���8����.��N�-�V��M���5`2
���	Wlp�_��^�d�k	4�n��F����S
�#��r}��)��ȫ��nM�u1����DD��3 ��cl�7��	��nADD�s!GIJ� �*)儩���>k6��GnpW7�p�wiS�����Ť���u���d2)nT�:uʡj����=�J<��2��hB|�U/x�ۥ�=�b$��ԔC�x�����(i3�{4STip��굮dR�VF��ڪ*�3U�>R���D;�t��"M5a�;����Sأ	{��� w�]���2�wk�a�	&D^%-K))48��A�H�vlp�O0D4U��w{e�Y���~���|Dfg����~��+UC�7��E/�GｗMD&����|ի�.�h�������(��Qh4���4)���n��j���H�ipժz��A��BJ�׀�d��ؑ�w�q��	�j����܉�<�����E��^mp�x������&Z����L�t������
Y'���w�e*�i��y��@�pXq���Mu�Nڌn���6'��+��J0áj�����PP�+++���UD����e/Ǉ>|�:�&����������׼��R�ƖiX^^R�35�S%iw66����,��&�N����hpR�{<�����V���j����,��|>D"��I�v����^8����+�h��Tz�k�3np��Ek���}�s�.�����wk�C"��R���&�$m�'����L����I�����U3�2u�{��N��躎��)�=Ţ�i�v�P�7M�f%"/;r�������c��$��|�����_�U�K![KK��A��aff����CzWJ$� ^�,5�3��.�fS�Шi��>I��Ba�I�4�~��VK�D�!�8V�^a�&�]6�[a�=# � ��cf/6����nADD�'%�s��܉v&5�K��ip����FCvH$���[[Lo���-���p�録9�4M�JV������J�SO�,���_���r#�<B�4�x�Mx��׻]
�X�t:b���ݓv�Z����Lq���&�D�)|4i�+�`��]��\i-��h��Z�="�j���nE:�ȩ�DD�� ���.b{m�� ���.�����z��u��
��-�K Kr�;��"M��A�H�u[��`�P(,~��T��n�\N�lQ�T�c�iw���t��v�������w�.4Ms�"r��׿7��N�� K������pD��E�abcC} Xz��t:1@#�J;T��ּ��ni-��T���!�(�[��QM?�@�	�DD�#^���.bP{��]�_��	��hb�ܣ�jLF&ڑ���l2��.Lpwܝ#5\4u.��lj*��.%A���̨4{���u��!�;n��ln%�7^wn��f�Y��R��V���gffΡj�ecC��=�����;T�7H)�<�a9��mv�&���l������0��h'��/�wT�0������] �]� �R��� x��E�3��@)���LF&ڑ�n"-�`4M�jL˷C(V�o����6J�՛�Lo�W2�ǧ���~���P�V޳�����[x�u׹]���G��ƛnr��1cbuuEyG>�C p��(�������5M��Ԕ�M>im@Z[��U��P�h4�6�^_��
�#���Y�ANpg�;�N<cM�4�{6iyN�����Ǿ�g\�=nADDΑ^��w�$�iy��i�D��{��n�h4M�~��t:�v��a�dR��^��لj�tZ=F\Ji��d�9��Z�&�@��
�i�`ee١j���7��-xӛ��� �1r�G������2�����rb��阞�q�"o0�rIyO6�w�o�^��Y�B�D"�4�z���.����h0�~ͦ��f0�=kpg#*яk��礢
J��ND�QWx��EH�B�{�� Կm���S�\(���8�u����DĦ�^��`E�+WB�qʄm�M:iT3.i�&�m65�U^/���[fff�׫�*��D?�W~�Z��lb%�g{�[ނ���&�� �v��P��]�v�XTO����bS���ݮ@�L��f�Ik_���"M��քi0ݮz�O�u��ꉇD^�w�`��DD�����v*{���\�vDD�,�%�I֘�N�3it'���#=���\"�T^��R�j���R���Z��f6
�����ƆC�xG8֗����h���տ��n���2�h���o݀7�گ�]��XYQ���bl��RiC��������t ^z��Ik_�ٶ�t؝�v�i6�w~�D?���r�����NDD��v�x��B��{��� ��vDD4~�xc���D;�D�w�����}�*6��'�J+�on2��N�̔�z��A�Ɵo�MO�(���}���9T�x{�+^��~���pED����w�G��]�X(7��v��H�Iix�nժ:�zjJ�F����T^g��}���)\���#��Ha>D^�騿gzY 0�}�DD�K ��vVƹ�=
�> �%""� U���&��	�Ή�ԛR�&����[^7�>n�H^��7�i8�lVy�Tbz�(H�D��k���UC4�^�������v��8/�Ѹ�4�y�{���n�B�:�4������P���(�K��lp�����������[[[���p8�@���v�BK�5a܉v��i�]��b�;	np��E�d�wanp��E�x�D"n�0�lp'ڑ��+�����B�ih4�V4��˵ZM<0F��������i��i���RIݜA�K&S�w�����!_?}���λ����.����χ;�x?���J�K!r���2"�Q���CD�M�6�t�h�Z�{R)������Lq�G��D�߳����s��R��4��ȫ��nMjp�^���	ư�|�
z�� ��vDD��0,���a6(0��hgLpwF<��0��0M�g<Nڜ���r��ɷ��n� �n��n3�.�DR92�4M��e+���i��V��J�9���<�,�}��8֙�v���㮻?���;��R�\U����Ki�ok�&4}i<X`3iқ4)�'�����>��;g�����Lp'�ܭI��NDD ~
���]ď�w?�O��.����!��e2��4&�ȋ���r�a��j�9��&�Q��ܷ��U2�R)��3���555��^�V��u��4MG>_P޳��
��]�\���q$�L�$�݋�b���>���Y�K!r�������s��^&�e�$,�]��#�Hk48������R���vc��C�L�V����;�����|>�2@��DD�? ���"~�86�߈�w""�(����jLp'z69��	6��C���3�����	��n6�;Kj�(�6��;��)1�ZjB"�d�p�|�#���s�"� �B���q�ɒ����*�ht]G.�s�"o(���,T��h8�ZA"�����V��#�<�w�}����4�l6��p���ٺ]6��H)�R�yB��n�����\ 7�]�����vy:�h��i�'.U7��jl��C$Q�m���gn���4M��Ǝ�����yK��4�BaFy}k��F��P5D�E�u|�ą^�v)D4A�>�l|����NO4�:�6*����i�wT���������16�ڥ^����Y^�u���Mj�LS�v
��hrI�9��a��ýR�g��Z0�w""�� ���E|�85�k > �v!DD4�"\���dd���	�lڳ��Y�������7@��s*��t]}�����n����v����L���|>d�Y�=���UC4~~���◼��2�h]u�Ux�{oq�"�H���؄C��~�Rd2�Z4ժ:Y<�TO����!��Hki4�s�D"l�����w�g�v��)A^�w""�G ��.��� �t�""\���;������PHL�t�V4��q���di�ys��EsI���xx�^�l�n�<d�&�����h|=z�^{��2�h��浯������2�\Q,����+�А����+J%�D��C�di�[*�w�Hka�Z���)�5MC$q����l2��h7�]��[	n�@DD{�,���]0>�I �vDD�7p��Z�M�D;�F�J��4��;'S�L���>�f��YM�I��a R3/�/(���%��%O���/�o��w�.��<��w�W��n�A�~�������*Oz�J&�����z̀	�����ki48),�{x��?g�L�����NDDC��s�.b\�o�v�?����pq�J�M�DϢi:B����Fӱz&8GJ��D��	�lp�K$A8V�S.���N>�_Lh\[cz;y���>��?bs9B�u��~ n�B�8iRP:�B0�ZӡammU���,�k�Φkmm����A�=�#�=�bLp�K��^wd�=��p8M���h�`���@ �v	DD�����v���~���]��?X����()z��6C5�%���e�ߏP�z��4M6��$
!�^�5M[[U+�l�tFy�^����:T�7�r9��Ґab�&Ѥ	�B�Ї?,� "�S2�ć>|��ۥ9�T*)���|ޱz��4MT*�=�z���׉Dҡj&[�����Ѩ���'��FRe�~��N�my]�4!؇ț��nMJp�B��ȓ^�Un��[��lw�P�<�B!��)4�<J�,���A��dz�]��6��CJ�j6�<�ai��^����gm���\.;T�w����rYj8"�<�~���.p�"�s�=��v��e9j��lp�_��~����h8���D"�P%�����V73Y�ҔN)��l���y8����b��DD�K���1���\����ƌ���j�hH"/�y[-�"1NNp�3���]J���I��Lo���(��p�~?2u���ښC���׽�u��׼��2���^�����_v�"G����s�Ri�3��n�H$��1��.lpw��&����R�	���j��y"�~$�qLp������L��NDDx�[���I �w��'"�1$��������`5я�Ջ�Lp����S�D5M���Mb1�f\�΃v����n�X,�`0hy�4Mln���N�lN��{;Ms������^�o���2��p�M7�ҟ�I�� rL�T��r9���z��l��4�t���&��֖���ڃ�L1NZ��"�`Z��r����W����p&�=�դwM�w""��M �����~��|""ڃ��n��n��Woyܝ!��m6�L���W�1��.r��z���N���k�-�酆����K�~�$��f�����	��Ƃ���?�G�f��K�`��Ţ�\N�ݕ�' ���hp�zC�����r��Қ�4��l2��	R`܉���e��J �^�b�;Y� x��[�� �ͥ?���Ƙ��f��%iA�ȫ��1ҘO��i!���Ai$�����H~��Hv�0�����w�a�ee����""#2"/PEQEQRW
�Ku�*�)@���R-# %�fF�[�n��������Kk��c��Ӵ>*ڎ��x�KB�P��qn{�8�d�����'��k�}���<�(u"#�g=;v��o��#+<q���}j4�:z�=�_�����+I��>�'<�> ���/֏��'\��a={�����&1����O����tqGQ֜����z�f(��jγ��>��G�ш�tp �m�n���
���$�� �F�l;ۄG�Y\tO�v�tp����aiiI�f3���`���X��[[��J�M�#G֜_q���@�̇cǎ��Ⱦ��F#=��c+�y��ߠ��c� ���;���]�ɓ'�'6%I�cǎ�h�Y�X+++l*��:�:A����h4e~�n���,�hvYw����������~������ P@�q�;��gJzC� 0���ɴCw�<�v�فy8r\�'V��S&�XY�{{(�ⲵ8��VV��jeO���H���+�}Ǐ?���ɓ'5U�s�UW�?� ����>�뮻.v@��4Չ���{��������ޞ�k�9���G�=�4M����
]�}��{{{{榍f3{��W��,� �X�C��1�?�� � �>d�&�ydu0�:� ?��;�(�������bup���T��[[s�&666	[{�$��ww�|챯������'���~  &�U�'_����:��;u��s�]�mn��VV+I�@��6knly��v��=W����:��xN�5p��nwb�  ����q7� B�_,����& �F�4u~�H�=S�KP8��vݓ��'Is3w?�����v�Jf[�$fG/:��������ԩ��*���kF����;��{��=tEPW^u����]P�'sv�m4�:z�h��f������~WC~�nW�~vخ�h���:ݐ�~t�;�����5�lJ��j�c�������,tp x�\I�
����74N� p`t"����e��@w?��hd�Z�z=���.������|Zv.�6�yd�&���U2���9?���d3��n׃ozS�2  �7��z��1v@��á�Q�z��t���㽲�B@գ�-�F�Ç�d�Ysc������hdtO8��k��~����=�p�� pڇ$�52��I��� j��Ҵ���1����X������
]ӽݏ$����k�E��4�>,..jaa!��4Mͣ�1��Ǐ;?�{;f���>��97�@�$I��؏��̳�E���$�)�3���:7�&I�ÇWV4۬��k?�����G|��|�L�����F�|��,� �\#��!��P+9mI��o j����$��d��Y�s��������^XB>KKK΅�^oO�!��}���}Y[swo�����:��%����}��;f����=�Kb� S;v�~��,�`�YϢ�v��g���w6�gܗ�WU2��'If���7�#?�Ta�����0�����'��%I�	=� S�$��r*�������  5eu߱���l4ioo/v@�X��l�ÚDg�����)ߟ�e�Xom���F~�������@�̇c���ۻ�.��0��z������4v p`���"�sｱ� J���'8;v,P5�a}�p��ِ�p_����;��7~#kΗ�Vw�N��6:���ΉI ��.���e�#!�mI?�� Ԝp��C&k��GI�ha��a��?������w��i[[�Ei䷶v����Mӱ�@�=F�v̮��e}��] ��?�~��������N��/���*!'O��v�'�5�M:^{b�ݍ��p�z�!�F���~�~�N��w �7?(�S�?"��fѽ ������D��,]B��y�����=�F���.k��:F�pcqqQ�V+���p�n�M>�Z-󺶺	"�F�an(8q�@� ����	�\� (������ñ� Js��	��V�]���\����h4����l�h{�}"��
c��ð�|Y��c8����F�ā    IDAT�h4����E�\tq��Z�  `J�Kz}��@�����/��  ̉�&òt	�籎@%t�5ք��XZ"��ʊ�{����$������fnD���X�l;z����i��pȆ̬g>�Yz�k_� ��կ~@��zk�2�Rlnn���9�"ѱcG��3��4��������@�̾�-w��:Q�Xsd�����uvH^XXp�C ?��;�? ����gi��� ��$��{��7��I���� �����̚���U�е�BE���p�}�2�;�o�d�Y��V�5�g�$��O�d>=z����S'9�3����C��
 3%I}�d�3���~���@��k�+wƛ�p�Ú#���i���s5&Hh\創��3!p>:�g��; ��+%��a�̕����+�� �a���;�p���H��ɇN��t�t���ZL���!�ÇW��oll�d>X!�'�!"����t�UW�. �{򓟬w<�P�2�RXϦ�͛t��ec�p_]%�i�:U����:7pw:�{-�N�\Zb]�k�ݚ��Q�O�=� %�!��E/3��VIO.�� ���pγ������ֽ�Z�@>�-;?��^F~�b2��9|���s:�����dWM���ʫ�������e @i��ַ�k��]�݉'��i���v�|�@~���㽸�Hʓqw�X7�tU-*MS�)��]�} x�լ�Z��`���Y�� (�u�^]�7.+�ޔ�=%}o ��r-ZH��"4Y���Ϛԥ۵V`��~XG'w��}h6�fg��-�1���СCΉ��hhݎ����;;;ܯ1�����0���j��?���.�n0�kss��5ǎT����q������ph6�XYq79@>V3k��X�kW�a�et:��碃{�V�=Wfe6  ��2�iY�WI��_ �T����&²H�G�=k����֢��X^^�����]�t~�ae�����b"ݣ#G�:??q�@� ��}�ݺ�;b� �{��{�7v�w�3�����lnn8??|x5P%�ok�}2���d9䳳��4O��������2���o0 ���f ���(�.�ߴ��;�� Ss��:����~m՟�%�GV��~X�VW*�c�L��k�Z�F~���p��@~I��ȑ#ί9q�D�j�0���}�� �}��>�M�9'O��QWWW�h4U3����tp�g{�
�����C�~XkS��ȇ�;0�~�F5Y\'�Jtp ��߰���ݒ�W�� ̱�1t"�Lj�Zj6�9����a��f��HAw?���T�ge�p��������oeeŹh��#����(��������e @0Ozғ���]������`R����]�}�/���9kn�X� b#��ܯu�'�����3��`��=[�$j6]��� �͒�����o	� 0�$q~���$X�^���h��R��%��B|h4�t:���i������4M�】��%���I����	��s��Q�����ER�n�?�w<�P�2  �w��!=��]�M��Z_?���Y�mmm�'��!���;w�����"�{�����dZ��Z�v��f��^��9�h`�k�$�v��� �jHz��o���^��{ �p��C&�H`Y�����X\���������8g�����e��'V���-�>:�l������ϩS'U��w��<% f�����n� Q�:E�=��hdv�ˏn��7�M���C�p�$�;yb�Q--1�>��ǹ���7�8����|de7  px��㾾����ʕ�  ���h̶G�8�5�K��kq�:��X�L؏v��v;{Rw4���+1�����$��ښ�k��P'�]w���U��] D��W�R7�pC�2 o�͘�V�I�I_���^T����qo&8t�P�Jf[�kwqGq���$����]ܳ�Z�h$� �BIz��o�3�~���z�~ �9b�$u��ɴktm �������1�aX��wvv8����Uw(bss#P%�ouu��-42ޘ)����9�y �u�FC��b�x����~���y�$:rĽ��Y�++tp�eg��^Z"��5gF������������;p>�s�k��$
 (�;%����g��;�(  ε��L&������au9���5�tp���fu�B~V(bk��5�9r������F�Q�j�r�t�M���c� ��|�ͺ�[b�xcuq��y�������/V���~Xsftp���H�8�������`@�=�u
� ]&�e>����{[�[=}/  �C�l{H��X���w^�au9b#��Ⱶ��|�$��[��w_�֎8??u�T�J��}���� �%�3��̋�����`����`m�'��5gFgq?vw�s��7��:�w:����K�,:� ���W��[$]��{ p:d�5&��yD�0�q���u\����|��v�Jf���!5�S�~�{�'I�huu��5V7L�.n��6�|�ͱ� ��x����;�3v�'O��YWVV�l6U3��4�����kVVVU3������ǚ3��ܐ��{���=?�5�8_�O�,� �H�UE�����C��  D�l{��!0��{w?�H��)�0���1����[[�0�>��P��t��l������% @�����XȳnwG�^/��$It��{c'��ɬ����NWi�f~�������%�����0g`ztp��lp �.������G��zIwy�> �9�̕��q����M��P����|4ѵ��$I�nw2?O�Թ �|:��sAs0h0�z.��h��vv��p��"���5���38P����g=;v P9O{��t��w�.�bcc���ښ���mo�O/���i:2�����`������7�M�<2����ǹ�j�aÃ^��4e~��t��&�{6:� y��B/]>�p�K�=  ��t�C��no��;�]���t:�n��^���Q�lr��СC��ywwϹP����	��b�|��PI�軾띱� ��z׻�C�	3a}��{(vw���7,-p�aw�ݰ��{C>{{�F'4���n(�Z*0i8$���
��� ��bI�\���<,��  Η$��#�L"������s�e�cuE����ʊ�8{+L����VH���s�n���e @e]}��zы^��0ks���s�2�6/--�Ѡ�;;;�����G��n���{C>V#&�~Xs�30���Z-��w �G�Q�/��A�j�� ��%�	�lijwl �M��g�z�}��͌�KKVw�>:�][��ȧ�n;��i�2֞,..:��i�jss#`E@9z��% @�=�����/joss�y�V�������gP5I-/����{tp���n��#+��8�Ne��h49� �=��<�_v�9b{s��Tٗ%}��������?_��=�G��$-IjJJ$��,���?I�T����
 �2���>;��s�Y<���#����}w��	���	]����>�~ggG��(P5�mm�ݽ}{{�F��[n�U�_���e @�]s�5������<v)���i���M9r$�kVW�8ʓ��m����677V4��]�!Xsg����{tp�32���l63��� ��i�'|D�,�WO��MI�:�)���Y������+$=YR�䚁X�������"��%=�����+�������g��R�g4��S�'j���I7Hz���[t�	P[I��y��B�8�0:���q��Zd���KK�CX^vܷ�	������ol��(ϛ����% @m��-o!�����Xw������/=��ٵ����Ǐg~nm^F>�\�x�"�D���n�=w��D_2���	^�A��N���j6��K��V��~���꾨q��L��>�q3\��.�t���k2OȎL̂�K����[$P�`����YI�I���������N��ؾ��"�fI�K���fT07��{�	�L=��y���sk���� k��ۥ���8p��
A�mџÇW�����
T	P��<�)��;b� �q�m���_����'c����{������w3k�2��������s��FC��
��C���:������6Às�Z-wd��p 3(����~O�<�H
��zt��zT�����mI7I�U����q�w�n��t���<�_<h��)���@h}I�-�7%����٫fK����>$�nI�Kz��'E����_Y���,`Y���>w�E	k��$I�q�L��#�����W��p�}ÓC����ooo�d�%IC������TP����mj4�� �Z��7}���������gإ�%�Z-�@�.�t-�}���v��:	�����qV)����<��S�'�:-[��y4�d���."p��X����~K�W�s���?:��i�ٽY�<�����4`j���]	�Gҥ��@C�wR�[�e���OT�p���H�w��K��?��w~fN�\xb���Љ8_��g�s�����,8G���4�V4���ܝ�����ߡC���[!
䳲��������@=?~\��M�� ������z�%��.8���o��>|8P5����:���6]�=����.^�h4��^�|p�$=��c?z=w��Z��p���,t���j��{��'Jz�����/d�q@��%=Wғ5�F��ƻ:�*{���Xp��P�G4���Gs�����Z�����wr�Wүj�K��6_Y�糺�X]N���u��Sq�&�>X���Q��gaa�9a>�oxb�z67�ގz{��H8 ��j���`^ԛ�,{��j�Jf[�����q~����X�6�M�ȇ�u�z���4{cL���.�S&�����}�Yw�I!PC�/�AI�%�L҇5n@[g_�8y���%����F��vLҋ��Ky�X���=�,#I��q��r���_�ZQyF�>&��wa��걃(��aB&A0�|�I�4M��3�UT��6��Y�8;��i>,..:?�ӵv����!V�p�T	����^����. j�5�}-�Qkֳ,w�]�!���s��ZG�y �Ԝ���xq��=��Y	��#����������J�K�G4��>��?IK�L�k4��T���	��Z��Q��~F�H߬q�{�������8��vI��<Lze�p&��mgGk���k�M>��=���M�X�+<���P�Qg/��u�ȑ�e @m�����xe�2��;����:��a�G��k��~�zt�/[��ΰn��P��
XP}ܳ�Z�/0��V�%]!�=���EOҿҸ��M����*^�q���p���������+%}��O�-'�=I����i����� ���ܳ�����:���(��{�8�ztp���aX�+<�|��9�tpG�=�b�  �������67���ٍ���	�0�]��;=�|���^�A��0z=�G�S��	��0v	�Ew̨/Jz���%}@҉����'��8S���8��-Jz�4aڀ�E� �0������8�����TN*�74�}�����-�Ñz�zƑ����6������`-FX�z�	°��nj���o�d����8O2���csj�����?-v P{W_}����g�.8��hh�;���k�	�����kn�h4ү���=k��q��Z�i0i8�iq�1_��ݒ����J��ݤOKz��gH����{�5��Ӿ�$~�!�ߑt����x��5>^�:I����<��$�;L�d!�L�����ݏ�q_&x퇵��q..Icq-���'tp�
�нu��׾6v	 03x5]�Q_�3���J�Jf��NW�����"�k�45�w���`�3�Y���;k}>Xk�)�����{�f������"�ZI�T��n�����n��G�k���OR�]���<�jʯ���wm�-��#�R7=I?�q��#�k
�8�lt�&Y�I�⇵�8�A��-..ݮ{�8���f��\,N�T�.��}X^^v~��E��������䥱� ��񒗾�0j��{��P���y�DKK�ѐ�ur�u�ltpÚ&��=ά��ܳXܭ&�@����*�]��#�R7,�vIo���ȵ`��to�/�&��8I/����RI?#�I�G�Z��˒�����qK.����qz�����$tp�ú/���{#����xB�~X�ۻ�.��Xa���:��� �KKKz	�PS[[[�ϗ�	��b��u�{�-��v��k67���=ﰰ��l��|�,�=ά����=�p*�+��$���[�Z�l$��4�~�3r=0��"�Np�$�'A%�6I�)��w~Wҳ%�#�I��h4x�r �L"��\�v��<����Y����E�Xw+4�|�$��������:v	 0s^���K d{{K�u���%5�,g�������z�C>v��@�̮4��˞�L���V���~�� ��p8�]Be��5��5����؅̐�g4��7�k��x�rfѧ	�3ۉ>"鹒�(v!3jG��H�G�#�k���rđ���>/��9��t��q.�u4����}��ww�]Ԑ��m�
M ���%5ً���{j��+�Գ����e ��y�ӟ��^}�2���C�㵵����	��@�=�}ؚ��͵�@�:��>Xsשׂ����-I�|2P1�$�N�[4dÿ� ��~!v!��%ݙ��܏Kz�A�r���;3�D��|�#�Y�~=v!���DL����X]`�,���G�=k�	��aܻ]:����������xM� `f}뫾5v	�����g#����F�ڏ�]�O�C�ڇ^��{���܁�r��je�i��
����&�c26$�����ȵ`��"����LO�(�K�Iҿ�]ȜyLҫ$=,�s�M�$��;Lxe�C2p>;x��MQ�#{�O�J�T��E-,���E9�co$ ����;�nu�C>++���h���] ̬���<����mw�$���؝���z�ǚ{ x����EY�F���H L��{6�˨���J�Oҗ"�2o~A�s%}"v!�i^�/-P���O�b�:��OI�[���.�:d�!8�u��uL*l��r��$6��a]�tp��N�a,-������1����袋.�] ̬cǎ���=/v�Ԭg[������)MG��w:5�����z���N�l�5�c��!����1�7Ҕ)�p�mH�VI�8��>-�I��̬�%]o}Q��{K�=��&%�S҃�H3����n������^����F�8W�V��,N��(�K>c���0�c����][T��tv�J��4�,//;?��\Ut��/�] ̼���ԏu:��l�|�4��{����[��Ύ�I������N�|���\�ō��]�bXW�E�llVDE}F�s$��؅@[�^'��z �E��	��&�H�Z��ۖ�JI�,v!��EI�K����k��ê�gL��n97����:��Z�@>�F�ŵ�m5ٯ��~_��EYG����:;�!�f�����`I���Q;�fS/zѽ�� �������j���:�J�V��Ќ|vw�=��w>�C��|��C�NP噣���n�I�p6��lͦ;6HwD�Gg�>�|]*��$= ��?s(O�����+�����mi����c��avpo1ٕ�O��`w�g�:��a-�q=G��0�n~��n�Jf���!�绻�l�@�<��u���b� 3ouuU��rK�2�����8??t����|vw��l���ȏ�{��fVS�c�Y2�~Xs�l$ &̋f��;*�_I�FI_�].��$�X��؅`�<_�󅗀;B���J��؅��/�m��a�B Itp D
L"x������b�\��8lu�B>vw�=�`�w��PE��ϔ$ �r�\��Ύ��"�~t��w��%:��`�9��8�a0�aX�ܢy0��ٚMw����$�^]���ɇ    IDAT��%�!�K���X��ԆLV��I��V���%�)���@>���J��؅ Lve���5��1�A���ȏ�a0�����������|쀻;�TM���_xO�2 `n�{Ͻ�ff�j���à�{��sii��kQ>XM9x���Z�y0i8$����p��4�w'���,�M�X̯�OJ�[�#��̸���p�$�c����8���b������.�I�l�>���~�����v���E5g׌�p��h���d-p����guD>Vx�ۥ�;���[o����c� s���n���,	�;����f��e�څ|�S�������5�$i��������#30oXO�f���� ����'��z���狐;�x��C+�ι�(�QI��Z�}@�;E�ɮLt�&p����qo*��v�1�� ��v������N����{�� ��s��YP9tp�ڔ��Dw�9�:�C��|����k��:��7tp��j����]�5�����A�=K�EY���/B࠾"酒>��	�n1����.0�
�3������{Q֑�l"��
�[�Ӑ�5��q��#��w̖��z~� `��u�]t�C�t�;J�4��~�<t��$�p���V���l�s���Z�4`�h��`�F��;�����K�~�C|F���'b�ZK$}cև���3$�^�Ŏ��k|$�/��NI��̟V�I�,�H�IV�6��Aw��1�a���|�V�yo���gqq�y�l����r�UW�O|b�2 `�<��׵�^� �4M���tq��ژL��8�aXM#_g�����p�3�b�PYͦ+6��$�U?����%ݯqV8�۳>p�����B0F��M���x5��I�9v!�/-:�g"L�&m�����c�ð��&�^�°B;toG��u'S� �w��`*ֳ���R�Jf�u����F��s���hX���.N���yK6�A��ܳ������Ib�~����o�ppwd}@�ex�����+��>�̏6�3�������4Mg��{=:��$��Z�F\�X!+$�|ݡ�n��;�宻���X�d�j�z�]\\T�l���3�>��`��E�._��4fI����n�E�܁i��=��%�X�z�BP�_�􃱋@m=C��}���*�D��G$�O��@��N��%m�.�!MS��tp�6��/0����&}ak6�J�$�s��:����D`u�B>tp�
�t��@� �---�ƛn�] ̭o�Q�_p-	����]��tp��zw�ޱ���Р�a��({���}����-�(k��M��~tp�Fw�+�U������%���E����n��Y��J���r0��T�w�.A�����.�.��,L�&m��)�c&	} �^>k�{=�؇N��{Vh�
� Ur�-�*��Z���w�ג�J��uo椃�vw���x��0�.^>k�1&�N��wVw�Y!0�wJ�b� ����.�t���c�o*ΡĴ��qWoZ�͏_�� �0�8������:��֑�t/�1��a,.Zw^�Qw�Ŕ$ �v����N+����O�G�=k.ˀ�1���κ_Q�10��h��ʢ�;�I?�ӕ�S�A�pG����E ��%�Y�"Po�]�I�����B��!;��sp/c�u�4�ŋ�ƘMd~X!+$�|����.�Q�* ���dy�����#]\\P���J	�à�x��1�拐�5Gl�
w`:�шu�<+#�OJzw�"�g%�-v��[%�� K�>���_�]�ؓ�zѹ%a�p6B����I[� ,�c�M>�Z���fu���������n�����pȉ��K/�T�]vY�2 `�=�Kt���.�%MG��ل��� �^>k���~�yx���Y���I��<��{6Wȝ�(hO��D�l^�kI�]jeY�3����-u��KK/��Ӓ��D�	I�]���R�L��F`�u��h4b�����o��;��;�(kQ�M~p/������]�Q7�xc�  �=�{2j�:�hi����`0p6�h6[�����t_E��0��Kƹ8�g���	V6���D? ��c���;I���s���-u�F��*i;v!��I���E`�0���p`���F��;x�8���4M����(L�����4��h�F��[a�J�}�M�K  �Ʀ#ԉ�����|��^>:��o<��=�h4�y`�]p��5o5�M��%	�Q�?��ӱ�@t��"��	�z����B��XMB^�����.��JzH�	xE�l��A`���q._��T�$��3�~���|ֱ�l"��
���uB� ��&6�Fvw�������w����ߓ��l�3���4^*�N�a�6kH�3p�4%����](���s���$�����]j��;�����]*�Ӓ~4v�W�O�;2�3�����Zk����̽�(6�a-
[�ʰu:�M����:V�E�*VVVt�UW�. p�S��Rkkk�� r��#�B�Gw���=���Ƙ�??������=w��G$}2v���Jz4v��$M<�^�풐ǻ%��]*�H�T�"Pf��ɗLV�`�
�Z|`��c�Fv���E�� �N��;f�3��,B P!I��Y�>�aPI�3��̌|�.^�q�=��ܚ�@>������8�!���
�[�������@�Kz_�"PK������-�$I+u���~5v���ƻ� /8d#�L���eS���{!��{q����`u=����f-�3�~������ Uýua=�������/MS����>I� �����Y�W��֚�5�̛�({ټ��;<�It8�����.�������R7,�4��.�Z`��{I�]fC�ɗL�!a]`?kC�B�h��٧p�/*I��p8�h�8eu������;f!J ���nd��@�=��ӡ���F�����k/�&�0�k�&b�$:�gk4�����)|L�o�.��j�9��ı���YM��#��K�"Py�_H��Db&:����l
��_so*�M��:�.�!$F�$e#j��l�g<#v �s<���ȌZ����f�I��:��A0�|�q��1���֚��Iܳq��'CI�]*�O4���8;�p�K_�����'$�r�"PLre#�L���0q�u_&\\��^f��#��ս��uq�N��=���+M�����+���� �9t�W�.ȅ.������p�)^���.ΚIQ����&�0�5:��X'̖$���/i�,��b,\���,���%�u�"P��`���j1����;0��.�ĕ��g-<0��q�A��Y!+�T�5�^� @�k��&v	@.��G�0_���u���c쇵�AGf`�@�q��CI?���g%}8v������-uHғ�����I�P�"P+�����.�� ��iH��@�=+|���_��1���gu����q�tz=� P]�\�&$ԃ��k=;�f��e��|���{��'����Z���@���ٸ_��K�T�"P+?�q�����������݁3~Q�b�����xS��5y��4 D
L x�\>�����:�t:��}�܋�:$Z�*O@uq���z���xq��@i�
���[a��$_G�=��0{y8I�/<��⭹|`�p�fܹgÐJ���E�v>/�c�J�`�����>�q�PK�����E���-�mD��@�0\���A��|�q�l"��rH���a�:$pG]\Kx *�{4���a���$!���� ����1��V6�(�7$�U�"PK?)ױ?�wW���#�� ��b�������t�4p�#�^�F�}Oq_��_3�E�%�|I�8�D�C�)�墬.�l"@����O|b�2  .��"=z4v��z�����8.Κ��#sq�ܚ57�|_��1��:a6�~�:��0�_H����@e��S���@���ƿ���1����p`���5��{���Y��j��e:�G��|�qtp�,���k� w�5��_D�ﻟ}�m:��@������|�5B����|؆�Iό10��v6kn��;8���ߋ]j�c�������S*O�P��I�]j��b�zjp�4"H
L�6��.�.�aX��l�B%c\�0���Y@h ��k������a�.��g���%�k>�j��5��8Q4v�@�}T���.�t�Ng��<�6$]�T��I"ၢ���n�"P?t�F��dM��3S�p��:��_
.��D@����������&� U�f$ԁuz�u����&����Y�Ĝ,����q.�k��hD�,�q@]I����Hҿ�]*iQғ���+N�G`�����]f�)I�&v���2	��1����;����k�|�b�`�e�1w:w�^����+��"v	  Ó�xr� �à�{����Y<;|M����M�1�_�pϒ$��Á���Y0����8�
��ji2����%}!v����ԚL�d$&�����)�.�ap-��ղ6k�.���&Z-WH'�4�¥�]� ���K/�]`J��n4j6�k.j8t���.�z_f��#	�Gw`:ܳ���������U�\ܟ�Tׯ�. 3���t"v�&_����dM��]�8:��A��|V�����Y�l"(��l:����ET^����pI�2  ��/��@%j�.�壻x���e6j��_c]����c0�4em%K�A�S���ߍ]f
U\�ewdJ���E`��%���E�^L�dp&�.��0�)��u�`CLqvw�EYc��3ƨ��.�X�N'v  C���%��!	�g�`�l�.�z�#|]��0�.�sQt�/cL�f �����5I,B�'�)\ȥ�ـ;gL�\�/�+��������^�D�6"|L |]>��c�C�$�g��k��1��%�|t��,���Kc�  ����XBB��w9��G��p�jn@0�8���1��tF#�Y�� �~���J���E�r&�G,�����L�I��E�>�D�F��dM�ґ�8{�	em"�:��1壃{��1��2 PlJB�.����1..MSg�Yk��Xs?�sq�\1�����1�ܳ�/�)�㱋�L"��s]&��?)b!��ߊ] fRW��vg��,0����61����1�:��!�8{c��#,	 ���$ԁ���JQ�&k#.�q�3�O�C>t�.����{rQ�:!5�Iiʼ:�cJ�ԋ]f�Gc�ʙ��N��="�����b�r�e*!G`�k�a��Bg��_��1ý��2�큵H�F��p�����; �ǥ�pG���ہ*�]t���峻��.�M�N|�:&��=M1%2_(�'$�M�"P)���ؐ�"i-r1��������>�D���p��dx���`?��\>�K>c\T�$�tto��.���9V����.�� ��Qvwq�~E�-8���cA����p��5
��ֳ�����S�0Ӹ��_"�I�L�\� ̴��t2v��E���l�/��Y�{�V~�]�|����⸎�`�F��pw���_� @NܳQv�V�Jf�Xe��;3����1�Z.�j�¦#?��Y�3X[�F$S�����]f��. ��Ćƭ܁�>� ̴��D��8+[��ΰ&^��A0�|�q�^���\>+�é��#G��. ��l���ё9����⸖���A#1 ?��]�W 7��(��u�!�h�*P)'%}*v�yܑ/��g��
~^|�ƙ�Rq���G��0��Y�tpG�5�M>|8v ��:�����e Nt�.��.g�"+�8ǵ\>�סX�� ��=S |��}Z���.�r�!�X�*P)�U��@��K�PI�$b���Yv�:P!3��{��z]>�86k��:ʛkU���F� j�.�:�[0]���70�>�Y�|\��#��5%�8g��up��!녲���$v��#�q�?�] ��_�. ���K6^$��^�@��|�q�^��F��1ƨ;B� P?ܻQutd._��ι	��~�Y�|��6U�=����F >p�@N����]��U�w�!�h�*P)�%}5v�>^��rβn����8ǵ\>+�`"��\>;��fT�ѣLG@�p�F���:W08I��=���l�(ױV�:P3���tXc
���S���\ ����pǹ�I �5�&^���e/8����\>:��/I܋�iJ��:��c�eT]��~�w���z����q.�����u��0�qT�Z㞌��x!�5�w�!�X�*P)��] ��L�Le#��e��2����%?��8�1E�%uw�.� P;tpG�Y��t���q.�=5��IQ���g]ǌ�/\��4���0���3�����謇��p�~'$��.s��@�Y]V`���a0�e�K~���k����.��6� @�9B��Fg�0�����G`�l��gϱ1�>�� ���@��] �ƶ���.�q�!�%����`�|.v�>&^.��0ɾU�3�����8� w�=`!3�
��%U���� ���w��g`k�(���ʘav�:P!3�9���C`#0n�F&9��BH\o8c�!i1v����] ���c ��O�IVà�u���_6��0��</��:�N�  SjwڱK ���A���X���8����`:�M�|>v�+��] *c�!�%����`�|%v�>&�.�wo`a�0�HP>~�E�q��qF����as��0e�s���1�峧%c?��ǽ9�m�0W��pF��;�{,v�+_�]  `V��q.���1����c?�'��I@��9	UG�0�.!�����1�q�Ü)p`������\!Ê3:ܱ7��)i/v ��#L����1�e㴇0g�!I �6'��^��F��X-cc�2 _�_�pR� v�+dXqF�!�%�q"v�;\ss� ����1�X>B���^�}�`�Qm�6ӑ P7lNB����a����\>Ƹ|���})3��~�����.�����2����vb��Ӎ] PO�|����8��`p���u\�3���a: ���s0�?���1.c\>�8��/�'ð� �2�8�M����. s�kNL� ȃPp�s|�qq\����c8� uGw �6'����n��q-G(�|�c��� A�b���5�3:ܱ7�F�8 K�$a0��#|]>�:f��#x����@�p�F�NW>���c��c���nǌ��/  ��'Dh�	qF�!�YI�я] ��������Bh�l,8����|�q0Ψ�v�~ P7tpG�+c\>Ƹ|i:r~��@g��_ ��G80��<!��!�z�F�0wZ�  �G#cVH�l�:`�܁ @��w����G3��W`VД yB�֌] ��!�v�,Z� 4�9 �t�	�q.w����#�C�ZF���LG@�p�F.cc\�q��0g`Z̙�� ��8c��H�,n�� � ��&X�q��1.c����H��#$	 ��뱔��s=��n�e#�c\�q��� �� ��8�G��qs@hl�  fυ��q.����Y���8P!3ξ�hT!I ��~�{7�������V���O���C`3L��k �	yB�F�g����@e��. s�h��:JLp�
�q.��:.�aBa#�� P?��nT�띎Wn?�\>���c��|\�a0� �@�"4�8����`��%��.q1�rPL�����8���u�q����d�UG` �N�@�1�݂�ǵ\>Ƹ|��c��2 ?�_�@���] ����    IDAT*�אD����!)]x��0K�$B�a0�!0�e#\>�^���=uGH ��I�>B~!��1.c\��0�qT `�-I:��2�8����+��/#���0K�$�^�ό�-�q.��u�/��=9�u���o ��I�:��Bh�l������u�|1 ��L!B"S�3�c�e��\yR�P}L"^G`��P�\6:2�����q�a]ˍ�j#� �ýU�$��s�>Z-���17�B�.e� ��B����3zI۱�@e\� ̕o�] ����lL��
�`p���\>6Ĕ��a�F#�獆;������. 0���n� �f�
���������]�|�q��Pg`�M�\� �2�8c�!�d�*P�Kj�.s�����x��8p��0_���\6��0\��3�����9wT���z�  S:u�T� '�����V�G��������c�_ �aj��������] �ʓc��8ِĬ$�hK�4v�W�. ���T6�a�Yt�����Z�M!��#I�p-{`wpg�:���I�m @�p�F�Y���&Q��F�򱉠|�q��08U����=9=%v�KZ�]*��;���`np����T6�a�Y����?_��M�cAv����E��1n6cT۩S�$�n��������gh��8�@`�l���@g��H L��?P�Sc��A���hHbE	�=#v�I��.5��K6^��}��`�2������=����:#2��1ƨ;� @�p�F��Y<�S>�\��G(�|t�f�e`�ƽ9� *��@�����&���q�p�e*[�p�������q-��Pp�b��������� ����:;x�~D>����{
s�E�Y#>֦�cA(�30�X.�{r:,�b��@v�� ��s=3v���\x���8p��� |]�4�����"�5�V7:��k�1F�� �{7��Pp��0جQ>�Z���`��x�F�@� �9nȍ�B�:�~�����~�KZ�]fޭ�@=��y�Dh	8˾U���{qV�kB��ٝ�c�_���=��&�5Pm;;;��ۋ]  ��p�����e N�;3���^�a]���lֵ��@g��9y�8�5�l�-���>��. 3oI4gƤ����s5$=/v�y��. �@��lIB08���!�-�|���g�1���S~��c����. �����`T^��r~>U2�^��F��!�|v�|��>��g��
�Y�
�%؇���\I��E�RN5$�]�*P9�BB�V%=-v��ErĄx�<�묉&�� �^>B��c�àS~��pN��� Up�ĉ�%  r:y���Q}�30��w9B�~0��c��gm��6��2��~�fa�Sx����E`��� TΗ��]*���`��!��r��=�0�,&^� �^>+Lw�⸎ðƙk��᐀;���_�R�  9}�KܳQ}�30a���,���gܹ��bAv�|�8��Bv� �Iω]fw�7���IIۑ�A��.�p�"0��] �	�lMx�ץiꜨ%H釵lu��Z<��xq�g���Z�~p-�o0p�1w�����s ���G�]`��{��wf��~���|�s-E�=��9Ό10�fX�8�Szq�0�%=?v�����;��K��בtw�"0��] �ɗl��I�4�D/��u��0F#+��DwQl�)��i6	����@}<�wT��L��8�]�����q�RhE�Y�|���I�t�g��S"󅲼@ҡ�E�R�(Ig�z��Ĺ���2|���b��1��)!�L \>Ƹ|VwqN#���.�8e��.^��i��D��#,	 ���$ԁ�L���v�MeK���#�5�F0�8kC�5w�u�Q8�l�1�%]�̤�b�ʙ�3;�s�Lg���W�. ��dm6�w�$���C��)}p]�IҠˈ��	����܋�Ǹ���K@}<ʦ$Ԁ��1�.�.�����a�3kS����|�10�F���,tpǔ��)v�9��YU`�G$���DIw�.3�5�@�0����.0��u��P0�%?��!�|V�����Ρ�;���/~1v	 ��ؔ�: |]>kc\��Y�5��c6k�uL'I���B��@�0s�+�)��@�|A"�7~!���%����/ٚ��	td.�uOf�� |]>k��uqtp/�1677���� �����ĉ�� L�6���]�	�e�I
�Ú_��a�K~�8��ܳ�F�1��%]����B�(p�۷J"y _^��"@nLpeK8����E��0��V��W�����qQi�::�F���:@�=��#t�C-�����~?P%����c��p7�H���Me5CaAq�� L������hIze�"03gT�s="��.b!���%��̌7�. �C7�lM����5?3E�Y<N#(�����EQ����+�c|�*x�Gb�  0<���P}�f�9/1ب��.G��8{�Y3)*Igȑ��\1����.��/����^�Y������`f�-���E��>+��Z��p!o�] f�풞��\��	������i壻x��M������;�����<��{�Y��x�����z�t�nw��=힞>}�mO{z!	p�`cll�l#06�$#H��$�U�5�`		��҂֪R�������2��{#��{c�~�ѡ�He�:NVdĽ�}n��|�Pȧ4	�{�?p�  ������now�wF2�������N����g{+�hp�.����=�B��t\�1�ܫ���?HzF�!0��e�]a�%^��S�4��������� ��h=��B:4�c8p �  Á��0Y�;�M��GHƺ������֡}���z�i��U8��2p:��q��pA�0��J���C`,}���ǩ�z�Q�Nr"���������d�thp�pNC�z�8D��w����=��t�c?Z-wH'��������&`���k5& �� |=z4�����ƾ�VI���0�("��1�s%-��I��C`,�ӂ$w$��ʡ����uI��db!1���_���,�s���ѳ�_��j�o}�Z��L���
4�c�=��C���
=  F��փ>z�d��"+L�zx�G�~�y�����ѳJ}8D �.�a+�ªhq���%�f�!0��y��q�o����p���C��T����C`rp��#���z� �>�^��\�%�������`���j�?ϙL�ϲ4�ct:=����  �x��	c"X�;�áH���A�zx֚����;�R>p=�c`0��q�cH��Ćv�I���C`l�p�I��B��� I�'�i����"���p:k���3~���L&��4���q:_�^�E�;�ý��$	 ���^�1hp�(rT�v;��{@���YϱU>�d����k��;����(g�&��ᙒ~%��8I�z������C�~5��(YI����Bb,�:X`�X�/,\�a-�s�`x���-�����<��a5��wL�X��q�k4&E�Xt>n}>��:D`}>A2��G/��%Ԣ(r��w:��}�։9D ����x���Ţ4��ϒ~"�[[�z��8���;�X}��k�-I�@ҳC��f}X�] G�t��A0x�h=�ϱv���a5���V�4����5��Pp��m4��a�)s���G�Z��9�q:�=����'�G���(�Er��ׅc�>I�<�7xK�T�;�!I�	=&B^ҫC���ip��5ZF�YC�x:_��F���t��>zVH��;&Ł{i�qu߁�B� $b��%�><�2�~=��q:�;{������@<y�$6ؐ���㡇�X���������HqL��I*�c��%=+��|4��#����t�|=z��G�m��9���r����a�t:�׌(���p��1<x0� �3;vL����I�Q��>@�l�.>,������G��x�x��a�v:V�Se2�ơ��<[��B���W�0�r۩�Ǚ��o��,I�z��=��(����pNg���w�����!���A:���wL��n�z�  g��׾z �B!�,�ZMZ)=�>�Y�x!�|�`�Y�>�튰���9�#���3����e���X��1�7IZ=��oJ���C`읶(I���*IO=��$�=���8��������z]&<<�ף�鴝��|^�L&ŉ��ՐX(�����p�6L��n���" @�n��&�u��zόd�;���d2����n�K)��:1���q� 4����=�U"�l�3��N�I�8�{I�8�_���I��eAқC����^zL�/���`�
N������v���9NG�i�9H��p;w ;>¤ ��됲u��|��Ӓ�
f_jX"Hw`04���v�	«ߖ���C`,�Q�J�!0��T=�_������S��|I�.�+���$���7��pNG(8���r�fX�&?�~�=k��ڸG24�cZ8p@�J%� �'��u�s�=�� )�����+��q��s�UD(xx��AS>0�("��jp�J�3%]!���q������C`"|����o��S��
���Iz���=&�纪�E�b-�`?8H0z�^W�n7��l6�L�5�a�=k��j�C2v����E��՝w�z �����g����P'��~��ℯ�E�{:��tpXL&C�=�kO
إ_af�OE�s��F_?�_p�0�W��B���,Io=��/������4��@�=4���j����<�
4[��K�rJ� û��B�  x��&c�X���zJ�L�R�}x�٤)X�䧃���ه(��!��gD6�ZtW���%�-��z���%�p�!01�ûߖ�oB������4zL�N�ÕW1���v���8<<���am>����G��=#��Q���<�z�p/��a`�p��q�m�����e��3Ö�d���^��|���c?�P0��aه8�1�L&�,Aa؎��x4�cDV$�_l�Ϻ!��C`b�%m��w���_�Ļ]$I�J��Ѓ ��H���C`rY�~i�Y� )p*;|M����^���]|�x���h��
w l[[[��b��(b����;�� �@���wl�K�V�����>�B��\�o6�)=��}��٬�3r?���aq�`��|�V�3�F��;F�%�"�fA�C���%����;�?&�ޑ��i�I��A���w`dhr����>8�u �v��Y��<�~�Z�F.Wk���c�>4��X$�>�^���)�wL�Z��o|��� ����oީJ�z �\.�\��v��^{`}��7#k��Zˀ��8V��Vó[�9D ���{<W��*+�D�O�A\&�B���ŝ�e�o�[G8���-N]͚�%]+NZaHf�{���8I��Y㴋�Z�u���G�~�9D��;xM�ݗz��HY.p�����7� f����^0�J%w{��^�X����Q(��>j�s�l���˹�g�ó[��Y�D�}g�^��x0jEI���7� HկK:/��8_��_p�Oo����@*��>(�B���b�+AR�t��GϺ��j�A2V�\�@�zXֆ���d��w?�����[�`���E� ��0I�Ü[[�}�>�Y����Uh@�zx4���Z#�֘a��L&���<����虒>�~���%�=��8]I��� w���t�=ς?�􋡇�l�p�e�` ��j~!|=<Z��A���Y�4��a��>X������}��=z �Y'O��]w�z 1�0�u�X�ip�����Ykj���a����7,;��s�*�e0w��%�Q�!0r�H������ ��q���lL�s$헴z�̅�~7���ii���F��n��̰z��:����l6K���G�C���Y��j�,��R�^��ӭ��X� H�-��B��\vܭàH�Xt�%����ѳk���Z��֗�-��`�ǳ>����.�t~�!02eI׉bd�����KҗF0fÏJ�����.����B���n��'��e8��鰞g��ó6�
��a��m��m>�W�>.#	�z+$�d�uw+��wL��o�9� 0�n�"���,�aN��(��{܇��f���N�C(�kݲ٤%X�\���Y�Z��D�8pF�2������E��Z�τ+vQҵc������ޣ�/'L����Qqp)c&!R�t���~�|=z�f�~X�s���yòBVs���k����2M;�(��r� �����[��d�s�jՔ&�nV��:���AK�������`o8]6K�M�n�58�./�ZI?zx�I�zL���/�=��-�	�Xҥ���?,�3�C���"L<�������"|=j"H��9lm.���v�?�Q�<{�n��62����r�����Нw�z �9w�u��?z �\.�<4��uip� ���N�u�ϱֺ���	�q:���fip�C��#��%}_�A���%�f�!0��t4�AW���Nx��w%�6���H�QҾЃ`6���#p�N��{��u��kӰ��q/�q�c?���b��>X��Rɽ��d�fJ��7_���C�  3��/|!��@��杏�ju�z񟭑L�Xt��l6��vS�h:ђ���G�Z�l6y�} �&����tx�`�.�Hzf�90��K�8��x�]��I��;f�Kzu�!�+ϒ��C�@,��+pNc�^d��}p�K4������j��<g26<��	^���Uw>^*�,�C�Vs>^.p�dٿ���# �̹��C� �:�i�GF2�g�z����В�׭���	���:�2 `����ۥ�A}���{�1y^.���T�u�]�_��'��z�$�,N�!�����k�݋0������]���ѳ6��MO$c��e�>X���7�<�����C� 3�������z` V��^'��C��>�mjF2��A������w`0��u:��H������H�;$�_�$S�t�����g���"I!^�&�O����]�X슗7�zf��hK���e�P����!������e$����|�T�)�+�c��q��Fgi ���7ps&��ܭ�|H�P �>j�lVQ�h����z)N4���a�����V�S�^�g]��u>��F��{$}^ҏ����?%��糒����#���6 �L��$Q�7�����!��Ѓ`6X���0������B�h6iO��<��<�f��{�6?�~T��1}��p�h ���|���# #��+�n�څdhp=�,��(?���&�6{a$�yNE�{<�1F��~���x�+Hz���<���t����y8կH�I����n��z�)M�bh�NC�u:��<�~�M����E�{:�u�����>4[�͈\.��4&�c�=�o}�[�� ��w��w��=0�(ʪ\v� ��G��>�L���G�*��Y�+�����30�("���;�̪��Hzn�A�͢��%=/� �:�����;B�I�J��Ѓ@���t��+%Q��Ң�!V��^�4�n׹ӿ��E�a�	xm��j3�Zz`�o�7
Ee2���R�Ɩ���X,rE�'V�gaa!�I n�o�w  �t��B� l~~^���w�? �No�)fJ�n�-�"�zZ�ۥ���,�fq?h���>G�ZZ���64�4�ǳ ����$�V�r��gK���zL�oJz���$/���'������_C2����啡�l�>�2��d`;�ף�l�_�	^�a����`��zΟ�L&�k��^O�����ϳ�����y�<7�.�Ӭ    IDAT��4 ���h%c�:����~o�d�٬�n4�B����l���-�鰚�eج�w �e�dd�t��1�2��Xҧ�ouG8�Q�?J��Ѓ`*%j�H�[|S��;0
�>"���?��t����K�ס��"�{�����5o�����vc��r�^{`�y�샵Ilm~"�z�
���������C���;B� S�[���y���c �7��#��G�l��o�u3�!x���t���zj�����7�!`;��u:��}���$}U�O�d�$���OIZ	<�ק�|Q�cj�b �WH���=Ȍ�$�\�͒�;�,��x�5��,��	�`�6s gx4���~�	��`]Yo�&��V�_w]� `j}���C� ��޶Z��4�t�#[����������/>�߳j��4{`�q��l���B�0��w`|���U�+��n��j���Qx\җ�|aҿ��K��F��$}Yү��Qz��/Hz�$�g{�^����u!0k^��Z$�ix4���ڼ�Y܏z�z���Ki��f�T��eEmE�<������ ����>�)�LV��u��X��x�懵��h�oEC2�Z����f��k����.�cM4N�p�f����?��IO<˴;_ҝ��U�A0�>��W�%�R�40js�.��yI?v��Iz�����e�Y��X�X��W(pN�l�N�u�)	��n����l���ש�+�h���^�9'��G��v��d2fG�JE7޸?� 0u����N���� V,���n��'��a7�p����+�k���=���8x���e2J?�c��[Iߖ�r������_%i)�,�K����e��.v��%�&镒H���$����%-������P$����tX��V[��6�hq�u�:�~�j��b��/,p�d��׆ ����T�ǫ�M�z�J�`�>��jՔ&�n��p=	��ʂ��f�t�<��f	����z�v��� �,��n�����L�H��$�+�Wς�qHҭI���;�ٜ�K%}K�<ˤZ��fI_��Ӂgv�e4ϲ"��i�;�k8H��gm[��H�^�;&�BQ��}�V��;�1�n��v��}�� ����#��k_�j�1�]���V���})�����03���	�+��+��c�V�����;eV~��3{���Xw��jo&�/��'|���w2�Q��t}\R�`���W��H�J�[I׋�WI��?au���$���X�ܛ,�Ĳ�"f��,N���S��~p=�o����z	������%&�G?���# �Ը��kh��Ĳ��ZL��>���th�� �"���z=mm�<�ZC�g�k���v�;	�S���
�[`�%���{$](����<S�5��,�g���A�x���$]7��>�'IwK�V���e\E�~Uҷ�?a�7�8��&��q
���4�
�>X�����y�v��v;�u#�"�yb5���p��R�8_XXP&3�R0>u��O ��N��O]}�1�][ZZr>n�'F2�g4���(�J���c�FC����"���b�}"ϳ���G̚l��8�v;��/�Jz�����A�8gKz�����G�"��<!��A��Aw5?6���=�K�e"������ �RVS�,#t��np���fD�@����Q��➆Z��|���[[ug#ZE���Oq"����5}��z �x���gu����c �R,�롽^O���}�nٲ>�!k�ak�}���ה,��A�tX{4����=^�C�S�$}@���gy��nI�����$����	I�+D�0h���O� �$���{%����;N0��^.�~I���� #�d�+w�t�5�4��A�:$H��Y\.���C�N�{Z�����Ŕ&���G>z �x�|��# �f���V��vi����t���Y�򑌵�B�������{�	0kr9��t:��I�c��ާ~�{9�8�����$=�~��O����vs/��v�� �I���n��I/V?�=����+$=��)��;0Z4��+nN��v��Q������h4ܛ�<�~lm���+�@�ݟJe�����RJ� �}�_՝w�z �XЗ���� vmq��^�z/���h�!f$S.�������y�l6�(�����-�z�'�{���mw���L�gIz���Hz����iW��\I���I�K���^I_�?�m���bG�L���AIWJ�7���F�K�+ԿI�5;a~@���U(�����t7�X'�u�]����sE<�4�^����ݛ�V�����rY�L&�i���&�n���G ��u��#���f���n3Brss���ip��Zs ���djh�l�ْl�'#�Zko�E��
�$�^�i�*�$ݩ~���K:+�D~e$����P�(�jI�t"`g����M��aI_���dA��>����$�kM扤��2���=,��$�xЉ��6֚F�o�YWk���r�f��������ZM����|��YhpOG��v�ʓ�D��{���n������37ިG}4� 0q�x�	���c CYX��4������:�^�<,�d�5k����4��`�6�s쇵�a� �(��?|3�:�1�~Z�{%����g�hw"���r���$�����Հ3.]�_l7wI��]�w@�Α�RI7I:&���7��/!�r����*�.�C�!�_j�_���
C�:k��EVK��r�d�w?���Ňg��Yׅ#�j��||~~!�I�[��t�vd2-,�\cru:}���Z��v�UW�բ���\.;o��v��g$c}6�ڪ;�#�rٽ��A?��3��óւ��d$cݚ�{=`�\���8V��r9I�Nҕ�ݿ"�����Ʒ@�i���~n���m��T�<w����n���U���?�Dj�dIү<����u��[$�&雒�R�'+�$���W��������^S�������Y��4��am�p Ǐz��X��e6������^�{�f�XPEl�{P�nju5�<baaAG�<��DӫR�8�'.--k}}=ŉ �>����e/}���B� �Z��ڏ^z`(�����77+�Lzb����Li��V(����N����bQQ�!�j��n�S�h:�w��|��{x� ����ı~���3$��Ϟ��bIuI_U?O�%IwJz$�ʒ~D���~���$}_�3 >����n����_�/�����$��'�y���7��'�;O��#��K�SᲤ}��K�3%=K������J�r���I{F�|>O�8C�8��?��;ϳV��u�5l�^O�Ɩ��hnn�|�U�sH��?�ʆ�:��Ǘ����)xV�Vu�5��E/~q�Q `"|��kU��=0��%w�}��qo��睏s�ޏ��9�㴷�a��YkoH��tX�2܈l�ˍksx�w FY��?��S��/���N�>�~�p7�����.~��y�gJ�~I?���r�ņ��v�sT�jp����'�����/���������J�����I��j|�-Ɗ���j9�Ug]�TR�V=06^������ro�XW,#�Z����,�	��`=�����٭p0	���*=�/0�h�Y��tt��W������n(��:|��c?��ܟ�k5�`��YkoH�Z&x����A`;��u:��# �dEҿz�lH:�~i�N�ߧ<�+,��'<Kd
1;����P�0���F�!�O� �b�� �����j�P(�e,�E��)���r�d��<�~����Z��={��>n��!�Z��<�X(���NكJeC�^W���װ��y�����ȑ#����F��˿z k7�p�<z`(O�u�y"�L�w�>X?�|^�\v��єL���y�Fl�TQ)�v^��n��3���`��.�?�7yK���� x����dQ&V�H{/p*����k��ڤC2֦1w?�ݮ�\[M�H���Rq�Nhq�4x���š p�t:���	=04�k�^�ؓr��l6�x�ݦ�ړr��{hpO���h���<��
�*���ݥ�i�>fe7  H�+��6�7���_J��=  0?$5ؠ�e-����u:x��Q��7���XhV�N�=-V���w_��ל�//p��{���u�uׅ �֧>u�|���c C�޻nl�������v�筀{5�I��p���;x�A�������t:4� �0t�ư�%}n�!  ����)p�V��n7�f>��JB��:���s�����t:mg3mE*
)N4��V4�U�mn�����)M2������JJ� �������V �A���{�C{;���྾N���V-�3��f��ͬ=�V?$S*�o?��%`�d2*��z=n�� ��:ú�nG�v|30��ǳ^/hp xp\�5�~ɞ+<| ��3ܹ&2V�w`�f�v�4�<��j�*��=0�f��\е7����Y_�p>^.�9 ��p��A}�c= ��O|��z��GC�-�"-..:��w��{�J���A�z}�Y��d�(R������Q��A8~���l���������@  WJ�����u�z�>  ��ba&V������K����tl���&*$c���������;177�L�[6|h�����?״�cZ����1_�,i�Z����C�x���켉��n�Zu��Er֡c��2����5
$S*��
^7�} x��g`p��u:� #Փ�>��Ǯq[�<|  b���X"@
��Z�-�{�p� �֕��2w� 0w?�͆�Z�(���0��D�m}��d��B����ѣ����o���q�����=�����������|��@p���w�g�Rk��Xk�����4x����ǣ� 0b7H���7�U�����' 02,��#@
lG�x:��T��~�������T*���)M2���֜�����4	0z�_~M� ���ῼ��c �X�Y��N�4��[\\r>^����tR�f��͹v[�𑌵f��E��k�۶���\.�=��"� ����F��ߑ�)O� �mX �G�؎�{:^���l�ڨ���T*�ǭP�;y������w"�Ɖ't��W� �����O<z��l6��%�X��,.��k����	��@�:��$ϳ܁����
��zܐ ص�n���|�%��� `�X�X��W"�l�lpO��tX�%Ӕ�u�7w67��V��5����wL�+.�\G�	= s��q]~�e�� �Y^^Q&���n�����,�����m\H&�ɘk9����=��y��6����a� ���{<� #�VI]_��g��fI_���  �'�qr�<Ё3���;xM���F�y�P((���������<��s���ֿ��yEQ6�i���⾲���$���j5���tp �]�x��	�b�X�UO�\�D��/4���\.+���[��Z�V�M�r�]VP������N�݇B�w`P�<�&q�m�{� �tD��>��π�$���� ��CW�YM$���s��`$�h4�������f	���뙇	h^�yv7���/�4�tk6��V�L&���k_��֜�������r�����;�= ���'?��c ^Y����s"�b��B��x�����f�M/��n�ʭ>$iʧY|xQ�Xt�vlm���*�!�l��QX�jp'� إwJ���p���G=O ��>$u:��r(���i6�f�u&�Iq�i�3oذ|��u55w?������S�d�ml��E��@$g�~�Œ��L�n��7]r	q f�%�\�N�z��\.g��ÜHnqq��x���,9@r����Mn��T*M�M���~�R�:{�fJ^;���D*⃺�^O�&?����٬����s�.�? �RU�徿����-I���= 3���Ԡ�=V� )p�^��V��x&�q�R!9�*�r�&|���	��Q����h��ڰ'��O��2�WW��4��o|�v���c @jn��F}��_	=����s���l�V����3X�B����a��YeH�*7�ڢ%߇~K�� ��!o�T���Q, ��%��MGq\�rI�Q �p��z�X4��YWrZWz"k��w?�M{�~X!`�e�U*�ǭ�@��Iw���=�1}.��-��	S �~�FCo��-�� �۳g��q�"�������䬵km��͹o�#��G��=��U^X{�^0��y�q�ݮ�f� �В��Q|�Q��$�#�� �G�{�����"��6)�M$cm�Y�vHfs�
�ϳ����77WV6�Ki��g�VVV��S������+�= ��_�Օz���C�xg�2d��`�w�.$���k��^�wO�e��`��r��k/��$��)�gm9�� ����GF�G�{y��戾7 `JY��:WƢ!������ڤ���kӭ\.����h��j�>E��ܚ�E��2�d��D��/'O�t��d�Y-//�8�����}z䑑���Xx�����W\z����3�w�ĉ���~������C`�n�е'z������	��a�����G�@�;0�\��8�v��D�; ``]I#�^rT�G%}`D� 0�X�W*��d-��,�ǖq��0��v[�f��L&�s퉵io]%��*�����v�Z__s~͞={S�H��V]�����z�G��x��ͨ�J{����777i��hi��٫R����'֚�u��#�����Z;F2ֺ/w`�|��{�V�w �W�J�kT�|��O�Q���   ��P#����A�����$����7k��T������;'���pi���I���|E���'B� �]�u��[B������ĉ�)M2��^��nH�ZS��$�L>�w�ݮ��|���9���<s� ؎�x�[l PG��G��2������� L�f���XVK0��E]�����t��aQ�P(�8�������ss�k���ՖF��?V�}qq��P=�B@ss����z�ޤ#G�� �9y���?=0�l�l?y�}x���o������a���j5n%� ��+���>n�#9k/���v�|��Ӭk�ym xs���G��2�.I"��M  ^�i �U*��g�u����0A�L`����\��������T���t:��g�Y�=��j����*-�N�JEo~�%��  o.y���Y�I����(�߾�t:�=*
��~d2�ϻ�n�C�Hƺ�^w��!+tM��/���H ��u�Ǭ�q �PG�F���:����)}  �F�{�L&�b�z`���m���g-i��Z@�-�k��ڼC2�jչ�[,�X����icc��5V� c���ݛ�$@���߯�}���� ���|������&������~Oz��	B7-/�?s�j5�=)�ˊ�l���vK�F#ŉ���Ff�H +t]����X,8~5�Mg�0�r9���X�� $�!I���u�]��(�� �pև%�h����=<��V	�����?����b5Za�
����Q6� &��_�:U��5 0�������ׅ����=���^��u���v���7�mnVS�d�Y{%����|ip��~��;Δ�d���B�1�Z��r0��;  �����K#�~��kS�s  ����n�զ-&�F`;k�j�A2���?�-gO.��VO�U�����K)M2���	��im����(������D@��9����m�� �]{�[ߪ�{,���,--��kO�8��4����e}fCrKK�k-���&��Z�%x퇵��A`;���\�L&�I  �%ݛ��F�]�^-��ҟ �`և�:b��s4$g��K%���P���9��O�n���,�C�Rq>�����$�occ�yȱP(rɣN�����ίٻw_J� a\s�Gt�M7� v뭷�C���c #u�Y����JE�F#�i�_EZXp��p��ZK��"�LE�:�us��Д���3�]�@�ݥ�($� H�)��i�ai��teJ��a    IDAT `�Y��X��5GC2����K��k�bn�,�E1���ژF2����tT����hq��رc������F��ůy��=z H�ĉz��W�c���{�������e1���%e2�[ŭV�<h�d2�����FJ�L���y�gZ�D$GS~:�=����yn�����\	 ֟Kz �?,���$�VG� Nv�;�8e��m���r�V`Z����!��*��)N4�� ��<�>lnV$�/�Je��������||yy5�IfC?���絴ġL7�� &s0����kb0��+��io�gnnN�l6��N�cސ�d��km�
�r���;�7nxb�al�o
l��}�V��|�� �ᤤ7���p?�~z �]�� ��v��.��X�^�&5����t>N���v��X��ݟ�whbe���`�ͦ66��g��n�����ޢ~���c �����n���c #w�Y���omm�Zu&�`VV܇���jHnqq��x���×>X������s?��-�H��è��7�T(���UV @o�t"�?0̀�$���Aw  ve�NA܁���͜�bQQ��[��dmZX�H��̷�aFr��x���Hnm���^.�U*q�O��x{�p�lx륗��{�= �z������%�@*�C�ǎq��OQii���n�Br�!�J�K�}��=V��U��d�(���z=5�4�g��=^�M� �kߑ����д�<�C�  �J��{��2M���z��y*�I?��{��(/���a#�"����ks�j_Cr�f�|Y^���'+T.���;`4�M��w��� ��f��W��w͛ɀiP(̰�uH�Y^^v�>t:B�%kp���V��w��;�~������U�<�qhp �U�R?]���]�� X�E�X�|����0�u�'���==�F��T�d��e�}�Y[;�||uu5�IfC�V3_���;;�i����>����z ���o�3�s�ݡ� R��Y�����zz̀��g�����&=�d"� 1�	�(��=�n�K�����.ꔂ;b�<^��v>��? @��H�6�"�ޔtq�? 0�M5�5t*���,��ݍ�4��a�y}�es�p�uُJe����X,�P(�8�t[[[s>n�/08���	�cv\}��ڿ�1 ��|�s������c �ٷo���'���le�}K���-,,8��[�7
y���^��j��xbܫ)M2ݬ�n���d2���f�  ��'�O�o�B�%�C�n�g Ƙ��H���\� )p&k��\��݇�����n��BA�\.ŉ�W��� ��ݏn�cܠ�ݟ~���@��~=z��x�<��	fF���k^������B� z衇��?�� fF�P����k�=��4�!��jqq��5�-[H�Z;�n�Cr���ϰVi�����EW�C�fqO��0� ��r9e2�7ͺV��|ܵ� �Y���Px��{O�oK��� c�ڼk�ۜ,v����
����G��3��9��}��	��bm2p���j��7hq��R�07������V��e/}�*�J�Q ̰Z���|��x-�L9��s$Ň���N�$l���ʊ3��j���I��/�a^���iW��}跷ǿ���[$=��\>_=�Xk��s  �"��C*�.I�K���> `LY�h~�7O�ئ^w���J4�b�][W�"�Z��<V,���k��ڤ�`��֜�p���1w���gp�ly����>�� ���zz����$0s����|�رc%=�>[Y7la04���*} ��k�#9k���� fQ��ވ�����; `���x�B�%�U�N� 0f�O,�ś��8��bb]��������5-�~X���%��0�~�"���JJ�̎#G�8/���T��s�M7�+.=��WW^�o�1�@��Ţ����_s���=+g�݇��\.����{=�w?2�Hss�u^n&��Z�����\����Z�� �A|[ҟ�"t����7� 0f�w��	�۴Z-����ǳ٬��b�M/����+��L���l
L�Q����֜��|��:�mnV�ۑ��������N�|�͡� 0C���Qo���H��^��n��I�AX&��ka����:|���8��;�-5����b��s�d��fS�ϵv�;	|(�J��l���{��U�n���.�� ��7%�y� t�]��%雡�  L�����vb�n����{z67�wB�~t�]mnZ-��A$�n�͟�={��4��1	�cu�]]�����z�&�q��A��+~[�N'�(@���ǎS���[]�#W��lp��G���5�����&�~�m��z����x��>H���P��=�  �F�M����#�ޖ�;��  L��X��;��ׄ�}��yJ���h>�L�j��\���lmVc0VS��={R�dvX�R���啔����ښ~�%/���F�Q L�j�����_׉'B���\.kii��5G�>��4���LEc�_֡x��Xe�m�H*�r���
��~p� ���5 �PM�E��xʸ�K>+���C  &C�E�XQ�U��^\f���k-�#�N��F��x&co� �ujnn�y-3���po6���׉ǝ�///+��������4O�s�9)M��x@/}�o�`$��^�[��{�'�(@�s���v���'�R�fv���q�ƟL&���E��XkH�*{��"�L�\r��Z-�Z�'�^$ v�P(�alY�Ͻ^/�I  c�bI��)�xx�$wm `&X�j�zJ�L&Z܁�hpO��\[�#�f��\���H�\�`����eZa<Z__W�ݎ}<�������D��jq߷�ln�����W��?|ի����%o��z�-�� ���G�Q��Mi�ٰ��h|~������⢢(��v��&t����0�U�d��]B����.�"�r��c�-  ���w��T�;y\�� ���Y�q�3��f�p�`�/�u��u�H�R�8_\t_��dZ���ރwz�����-�{��1�'�8�|<��i�޳R�?����{����c �"�]�^}��=���J���k�����Y�R�����_�����QzR.����c�v���8L��ݔ�A_�=��vѸY��x_ 3�)�BI�Ѓ�j��t���=  ,��S��p6{κy���m����X,*�����y��Ar�ʆ�q��
�Y-����}:q���={��4������p���s�9)M��w��]����B�`
�߿_�α*BRg�����2?�apV��ĉ)M2���3����+��<��K����\.���z]mmq�5p�|���K��np�w% ̼7I�V�!�4nwIz�$>� ���d2��iۈG�;�]��3|���)M3��w����}��4��e�K�7o��O<�||Ϟ�� a��z=��5�֗���У �`_�����?��� fZEڷ�l�����_6�3?�p��np'��u�����䬵��M�}�3��j�:�'��v��jp��q� Rt����3������C  ²�@ģ�ؙue'aI?�ժٖ���_�����ye�ٔ��nV���⢢��ڗF�af��ݿ#G�P�ۍ}<�ɘA$`ڵ�m��忥{�7�( &��߯���7�h4B��w�^�r�[��×ܞ=��5�v�m�3 �ry�h_��|{d�<p�#�ͪ\.9���;?��
k��U���m�  �t%](i,-�1�.Io���C  �!�{�܁��w�����vU���kZ��h6��pL&���ϵ�ZM�V����LFKK4��d5���Ii���n����s�97�i�񵱱�^�=���G0Ay�]p����z 8�=��ƺ�������	�<y�ГG������͊:�NJ�L����;�	|�������uu:���bV��ߓ����k6���%;� �j�����3�����$m� 0�h'��@pؑ��Q.�������k�*�f$g��[W�c0V�zee���x����y�?��/�c�=z ���ú���ȑ#�G�+
�mL���ƞ=�C��!c�
������������N��Z���D��Z�V7S�d����N�P=�ز� ��u���C�2�wI���׆ 0�j4�����*� ��np'��1?O[�/V�uE3��6���kfmm��fE���YMq��p��	�m�t�OKi`�>|X�;�|:t0�( �����u�/�@�s�}�������Q�����h�p��Z#�ؠQ�k�v��>Xk�ܼ�w`whp��l�� �YmIϓ4�o��9�.I�J�B�!  �Z�߯����lS3^7���\����p�5���c�Wx���jm��k��ݗ�4������wc�9眫(��$ ��/|��;z c������Ez��C����c����Yg��||ss�ГG�BѼ)r}}-�i����e��!9kM�ZF2�L�R�����v�LF�|>�c��r7��z�t��/��2�;�]I/��'O �1և(�ݬ�"�Y�n��W���K)N4��4���jp/����X��as��n��x6��@�gǏw>�w�^^KF�СC��s����;;�i����C�E^`�0[677u���o;�(��X]]U���>��(�`܏簞O��������s���܉���`5�p��\v�4u:�'&��n�w �in��'��Hb���I�z @�̀{��-�y����f��9�"=�i4�Ƶ(��&+$�n�U�ם_�����ݮ^\YYIi���YĿ����ZZr_���U��f �iOs7o���{��K^�bH�����D���7C������h��I�-N\�T2[�	������[��!�L&2��r$S*����b�t:�׷R�hz�͹��iovV(C�0�hp ��&�9�&�
�I�K��n=  =և�^�g�fق��̪z�
����j����QG��?�&�����4�Mml���V!v��!ws���
�3�3�y�z��G0�q�JE/��}��_=
0Vr���:k��k:H�f���l�p�u�����,,�+����VK[[��}H���k�v�������]�7\sK* ̘ߓto�!����{Oҋ%��' L�¤$U�,��Y��ؑ��NX����jWBr�F�uU3�[[[s>���l��`�&��{	��#O���8��j�f�]wݥ����9z lll�E^��n�-�(��9�s��J==�����%�g�c�ho��\.�T*9�f}ݽ���R�����r���k���/`g�B!�c���8�z	��L�{I�=� &i����牣� �'�Ro��;�#��!p������K���N��xEZZ����ر�������·N���G��s�=W��$-+�x������?O�
=
�;vL�?�<�y睡G��Ӟ�t��'N��eyr������_C��/�f�j��lP�`�Rn'��Z˥��܁ݡ�=��ރ�; ̌#���	�_O�N���z @:�SU!b����a؁��KHҟ����iJ��ƽX,���I�������k��l�V��^wN:�,Z�G�С��������ۗ�4�d��w����{�y��У H��C����K++���w��>�~��ٻw�s�����&&��v2�If�U2@��k-�ZFr��U��*�@�5���#  ��_.>q�<�p���$}9� ��h����d4gl�hk��n7��\.�b�}�0��V�f�:�ϧ8���v;����ɭ��7�	��g5
p�����g<�)ML����<G��w_�Q ��c�=���~�-@��?�����j����)M3[��J'NW��Mi�ٰ���|���?�\�l��T6R�f�e�Y���5��M��|(���f���w:5U��
��p{ @�%}&��1�����$�k�  S�
�̺��H`6�T��N8�C��5[���m���*��D��k3ziiѹ��?��/..��1"����������eǎ�_�|�s�ݡG0����{�У c�X,�!�Ç��(������5�abf~~^�B!��^�g�Gr�2��
����y�_�u?םN;���M�����yE�$���a�>t�U ��$�.��5�������C  F��0�����.�B0��E`B��X�=���"}��pܗ��bH�R�T�Պ}<��h��l}}�\�߷o_J�̖Ç�Ӊ��D���?~\��}��=
 ����/��=�p(`x�ӟ�L&>)�t����3K����<|���t���>Y7�mnn��&�U�`�A 9k�2*捛�y���Q~�Ɓ/ �iG$=G�{�o�Mj�]�>&��C  F�
��j5�}�;��9�uiqq)�I���i7??�\.��4Ӯg>�֦6e/��F���Ov~��g��|>��D�d��jz�KC���C���O~�z�_���F�Q����D:�ܧ9��������Ji�ٲo������N��le�].`���X�V���p)���npw� ��X��Av��� L����J:z�aLr�]�^!���C  F�
��z=�j����<4#;��==��;���?[[[j4��g2xdmJ[���Վ���LSψ<���Q3�������׿�z�%od��P�^O�~׻��?�CB�@g�}�
w��z��݉�H{��u~7P���d������s�����R�f�Yϵ��䬽	ko�U��5��# ��z���=İ&=�%�$= ����y�dgy&��侯��WwW��Z���c[� ��Y<�1��`;n��1�3cپ��q
�=6"��m��\`���nFx$$jaRKꥺ�%+�}=���@B�ߛY}�<�/������<��~�K��p��T1�?6�]�������p��L�+�J �_V��|p���a)�JJ���I���p����f�B#����V+��Ս��<!ЩS��я|�i�D�L���m�]|��&2Q�����y�VC.ǆ�QH$�p:US�t6�,�('��<������N��Hq�\��5�=`�RN�~�O��\f�;��x�lp��i����}�=]"���� ���E�7���_��"�	$�TI��v
��RJt�v[L�&V4�:��՚r/�G:(�D��n�J�"����'L��t��LF݀�JM�T��lm��5}>	uB$��}�}x����f�.��P,�k�z+������R��p8�HD=Elss�K�tp���|>�L��%�=�b��l.��D���y�B��
��?g���h�Z�4�z��u�[b�.�	����C6�M�g ��D����w ���Z]������=��5��J�#���I#j��n)�=�p��@R��t�M�K���ϣ�(�^u���~Z<Y\\2��������������K!"���U��_�y��K!:T����;�vwwL��^�I���t����&��r��h$)�A�#��I{���/.*�3���?&���h��z��h� ��z4�!2)� �' ���E���������J�
���(҈Z6��\.+���N'���f�ϙ�n�l6�v[�
&%��躎��-�X,��DCZ]]Żny'���/[]
]�?��x�-���ŋV�Bt��|>LM�������f
�($�I8����u]��>܍�v���-i��#M�(&���r�{���K���m�EtyN�.W��>v'M���"����� ���#MR�; �6�G�.����Sab�G�.�	����i]�Q,��R�.������x��LF�5b�+װ�}t������i����&UC49*�
>��㮻>���FD��u���n��o������^laaQ����iR5��JM+���y4�L�4R�{���V��R���F����x<}��Φk1��<ҙ܉.���j�TN""�(����"�6i�u � `� ф�n��ܨT	�����w�8P\�\V~�{<n@H�����(�j�r�C    IDAT�iD9/�V��G"Q�|>����f����=�Tj�?�x����~ ���"�V�P��~��q�]�@����ED/�t�0;;�\��fQ�0�d'��rM:��NOÓ~��v��%�)���%^5�����u^�0P0�>��Dk���z��"5�3���hb� �Q��w X�f U�!"�+'&6�M&�(��KtY�Z�n����ͦk�t�]����&�S(H��C@N/Ž?6�/�ˢ�n)�LM1�}T��ה�5M��S܉�G�-�|'��w�.�Ȗ�:{��x���.��К�����R���X7��I&p:�}���b1#�X��r��w@Ñ���1�4y�Z���i�T�d��|ʿ��N�Z�Ċ���5�lp'"����z�z��  ��"�	 ��ejAl%�<]�Q���C�Bꑠ48iT�tXB�+bb>ӕ�#RG"Q�����k�P�OOϘT��T*�r����9�����������ʿ�����.��V��^��=���:o��w�qA�f��tp���](�ϣ�R_���!���
�\δz� Q7�K�ip���4ِ'�E�d&�_��񼣿n����'�`ѡ��- &�qnR�� ~��"�������D�'�唨�JE�?d��Q��^�1N����n�R��L�4�:ɍ��N�)���aq�3����t:177oR5D���l��~�?��>��D#V�V��������z�fu9D�Z*5�W�`$M��s�\H&��5һ/�P��K�Z-N�5���F P�)�A48)��X���(�Y�t�AdgLp�OJogѡW� &z�e���N iuDDte���7��r8��/�]I�Blp7��U(��c16�E��$�x\}�M���rb� S�G'�ˊi�i���D4z_��񶷾g}��R�&����=�����ۿ������tD���l`o�֣�JM�����7+mbE��H$�ϥ�o4iO�^���|48&��G:���g����v�h�/ٱ����P� �e �bu!�f������� "��)qcGI�IdWR�4�W�T��v�>w�\���&V4�
�(f&�K:���ix���Ƀ333 �A?*R�����,/akk���p�]�@�ݶ�����vq�=����}VWW�.�h"$Iqess��o����̬�y6�/
�p\.�ڐ�fL��b1����'F��z}�x<}���Tq�B�I��Y]���V^�;^�""�h��^��0��ҷ ��q�!"��(��v�0��r����ύ1�躎rY��#%���yu�����I��^�����������|�����ߨ����P�,-e
�A:�>{������kkl�%��۽K#w�q=�t��Q��n����-����χhT��#�C������n3��`R���'F��D�{��rYhB�s:��^�4I�Ȯ�ޮ&���nR%DDd�;���E��.;E o��#"��$�\q�X-�w��j����M�ؔj �ZJ����ZM��C:��5�M��L"�4��(��V��5R�!������T����H��M����q���o��?�9�K!:�N�>�_|���跿mu)D%������ۼT2BһO��F&�oR5��L�����,���x�k���I�L�PHjp繜Qzg�/���uN�"���c��
܉�&�� �.�Lvip�u ���"�CFJ�h4h6�&Us�0���?�)5T�צ����\ҁ^,3�{����SSS&Ub/{{���T��8FhssS<`=z�(T��D4�J��߿�v|�w~��lT#D&���o?��~��(9��hG�S>�u��cS��3���t�I��4M��.M|��Ha�z�zݤj&_$�����TƑ� *���y�^�Kk�&܉�&�W|��>��v�{���6�!��	0-B��D�I����c�RI}��وj ��=g���2��u$���1����U�_w:]H&y�`T:����15�	D�p�}_�Ͽ�f�s�)6�)�>}oy����V�B4����~���æ��D�b����DËFcp�݊�x��#5��ry�*�|��!a��Y�a�g�w�~��ޟ��ʀ@�������7������c�� ~@��B��hp�K��lg>��MuD}H��(V\�ZE�����7�ip�|^���v{�KF(h���~�8���W��Q(�kff�I�te66���t�k�=fN1D6T*�p�w�}��\�x��r�����~�W�ȇ��1�hTz{��ukkk&UcO�;O�^G>�~o��I��
�"��,WO#��hp� g��N�
[-�"M6�e���^��%��F��<#b�;ѡ�=���my�юo4Vb�;ܕ�L�&�,��=�Tq
�wi�-��n��>R�N�uq�x2�2�{���$/��P������rM(F<�0�""{:��x�;ގ?����WD������{N�mo}���.�h�A�"o:�F�V5�"��4R�i嚽�]�lz�)�ia�̾I�؃����W����ni��P(*�&ip�C!)y�It9��q�W��P�ñ�����8� l{����:_�^ �1"":��a�;�e5uqD_02���V,�âQ6�IJ�����W4��}��u<���?��&��C����\�4LO3�}�66֕� ����^��ӟ�3��/�O>����Y��O���.�y��V�PK4jǎ�n�Y[[5��J&�p���5ҥ`^(�ϧN���h8�:��Z���d��Q�=Zi��
��M��f���D}x�>6i+4u�K "�+��& �~��s�; �-�_�>�%"���w��0��ΤϏp8lR%��PP~0��Xr�{���f��v�ߟv8L��v��LF��?77oR5��h4Ħ�h4��"��}�I��[p�mcr(�F�P��y���[����Ad�`0�TJ=�*��G�b��٦���S>/����3SS���j����B�=0����w�HgŢz"*��I���Njp�$"���F�����uX��� �� �2��ND4֤��R��<*l%�O���aJ��2���v#�X�d�����?o���	�v;���㰧��#��`����Ձ@�߅FlmmM����|ܤj�����K_�"���7�w߭�XDt�u:|��Ûn~#N�:�N�[�Df9v�8���5s��)��+^"���5�{I&���Lo7^,�Npg��q�~?<O�纮�<�@���r��^D���]�^WO`�;�XKx=���.d������o ��.���.O�	���5��OX�$#�3i��	���v���[�K��v;(�?oi�3'�I+�'I��@&��7�dC�2�z{{��p8�d2iRED �bw��	��-o��ӧ�.��P?����o���~;r96��)��ws�,�E&�������R׻�wt���C(�`���� �^�b��|^8@����2/H:{�e��|>��%�5&�Z{ ^�q�lp�!6��9�!�����Bp8�g��r�ώ`0 ��iR5�Oa��G�p�+i�3g?��ư��f��躎�]u�{*5��eRE���zI<�%}��VWW�я|����3�X]�y����[?�s��Y]�-;�,�Y]]5�;�0;��Ļ���V�eR=�!��7�6�LJo/�+�]7�>��K�q�\�����܉�a�{�N�v��7����ۿgu!��^�s`�;�ؒܹ�֏��@8�w��i�ZB���P�)�F�>���n,��=�1Q�@�VS�4#%��loo+�;�NLOO�T�=�j5�A(��Tʤ���G}����w�����tZ=u�h������;�����9���B�p��z*O6�A��4�QJ$�bS����I�؋�N��v�I���'U����\�̡��l�^���>4M�{؛���3!"���� �ou!��/�9 ��܉�Ǝ��Ub���F��+�I(ҨP�t�����xL�f��Et�ݾϝN'�>L:̖���`j���D#%ҕ른����K��!
�U��6����w��7��o��MX4���<��ӟ��o|��2���FoyY��s�ҥ�bsһM�^G.�KFs��b�o&��V���w6���r!P'�3h�8ҙ�ۉ��z�l�V��V�@DD�y���	�Glp���� 5�!"��9�S��D�I��9�8�V�ZU�&��Q�ݮx� O�T�=H��~��`Фj�EJq�D"�B&UcO�z;;��`0��i��Y��j����p���GwށL&cuID/P�T�ٻ��nz=>��?C�R��$"ۋFc��c&�/�Еq����靝m �9�H2�T6�u:��X`�p8����������pm��U�x��&�"�9HS"��L�dcwR����{"�� �* OZ]ȸb�{�� ߊ��Ƅ����5)]����e&��Ij��c�rY�si�<�Z��ZU_�H��M��^��=1Օ)�w��%������iܒ"�Z�N��nz=����F��V����w�7���;��J��1Xz��	�����,��ߥu]����6=�~��f3�'�P_�)���t8��(Ҟ���KÉD��NtP>�zڄ��2ѡq�k <cqc���j���ز�""��+�2:��I�>l%꯷Y��3���+ӂh8�a܍�ͪ�C�<�I�؃������v����U���A��5�lo��Q|>?��xـh�<�T|�M�����`�(��P(�/���u��w��	���������N�Q.�M�Ⱦ����l�MM#�r��Ǖk���{4<)�A���H{��"܍�v�����u1���Θ��w"�C��W�`u!㎧�����~��B���Nz��un����a8�N�� K�v�ZM�&b��Q�Ðp8���WF�T���v"�>����崙�� B��I�؋�X�r�x��kk��v�O�[���2�""T�P��>�I��U7��>��/Z]M����ѝw��׼���?��
�1�i� ��:VW/�Q��E�1A嚝fv���TJ9����"�ɘX��s�\�TM6���p�?�B��ӌ�D��+�*���஦:�4��DD��:��س��C��Yp���""��7��՟�i�՛fDv&���6�ip�j�V��sM���4�\N}�'%b�p��"�u��6Y�F�\?���L�ƾ��&677�k�n7���L�����l6�/~oy�/����CY]M�'�|���1���7�ԩS�c"������r���*�����]��l��zD�w�l6�N�mR5��H$�iZ��VK|����Ba��[��F�R5���&���w��?Mӄ	��l6��v�>W�m%""S|	�� ��m@lp����Յٙ���w5i�0���� b$)�]�K��f����А��N�S���>:;;���H���&X[[E���2 ,..���TD��������A���w���%&	ҁu�]|�����[?�w�������'�1�t:q�زr��wq�ҊIٗ����TJ�fgg���#�r��ǔk�i�M
c�9���(��Q��?o�Ha:��:���x�<�P��w��#"��) � �[]�a������ϭ.���.��w%6��'m3��X����=S�p�ٜ�7���F���~?B��I������,���k��X[[S�q:�8z��9�{�'��.�t��W����:������wߍ7�|3~�7���A.$nmmq
�	����$]��K�J��i��Ի���G O(�Ka4i/�PțT�=��Lp'���gz�J�ΞI"�1��� p�א��>�6���G ���BDD�`��Z4ʆQ�~J���������X�d�ܣѨr,.��i�#	��!�T*�MLq�N�������i��L���4�C���y�*""#����O��O�W�
���A�>}�)��"�n?�>����׼w��	���Z]��vciiI����`u���GM�4���)�d2Y^4��=����B��p�FG6�3��I�i�xv$M���|>垔�wQ��M���p���V�0֤wN�!"2]�� |�t �9�Ox3 vR�Hz��&�܉��v;�V+�5�S܍R*������������4��}u���4�GessC���p`vv֤j����ҥK�5��ay��9�������_������׭.�,������}7����~p��f0�at��2�N�r���*Z��I�W*5�W����iR5��v��ŕk��=���i��T*��@�pN����n��p)I{��r�.s�������w"���p����B36�_�p ��m""2����n�Q��T�,
�SDv&���DxI�(���)��� ����f�����&r�|~�B�83
�j��:�m~~���T�}���\V'�MM����D4ޞkj���o���گ���%��>M�J��{���_��e���e3"o�@ss��5�fC�XJƘ�_P>��j�;?��TJ����v�@�4e�?scI{��B�����J%^& Ra���4M��DD�y�Ox��B;v�]���� ��ŵق�iʗ�b��`0hbE���i�Ţ�d�Lt9�bA9�Y�J���s��X�?o#��%4�Mňg�D�����5�J�j��r�=�J�\V_������T&��|>$Id2�&VeG:.]�����e�UǏ_������v�x���������g��p��7�u�=��'L�^�7��0N�>����e�j5�K""]u�	�2�K+��ld�P($6C����=zR)��L&�s:]b�H.�F��`� ���δ|��<�T;k����d/,��+ � ou!������j ���,���h�9��Y!���,�����)Q<��p������y�;]$��˃B��rY����}�H$��n�tzG���|zz++M��>����h4���?���_`��	2������A(������L���F��l���������^/~�g~7�|3^�MV�G�h4���������}��Z�Z]�@29%�'W�U���T����/*�w�����-6�J��hx�x\y���n��@�C�P �����N'���r�tFAdgLoW�����fJDd�?� �V2)��n�6�� |�� IDDdn��E��L�W�ZE�Ղ���sM��Q(pS��r	�v.��_K4�w��T&�d�e�{<� ���oƑ�}>����������±c�}�$	6���ŋx��_��g��-//#��C��}?�I�h4~����?^��W�W�
7��*�R)��#���}<����<�����7�h�i�W]uB\w��N�1������:A|ww�vˤ��%��V6�u:d2ܳ2�t�&�����@�H����N��=+E"��J��D���HD��|lpWi4��DD4Re ��sV2i��n���; ����BD4���K6����3�(H&��>�F�lp7����������blp7P6����}R�n7"�0��T.�Q�Ք�2���<,���-=z����v~~�ϟ3�*{*�����U^�q�=8z�.\8obeDd�Z��ӧO���� ���%�x�x�kn�O��O��lJ��t:xꩧ��C��_����w8�F�d�\.�)H&������T����4�����Q>�d2��8R�{6�}B#IS
��</HJ���&����u6�Y��w ��ՅL"6���S ~����k!"��B��l޳;iÒ��
u���	M���sB�;/���n�T*!��]�LN���`R����G��l"�Ncz�c���VW/��b��]�xSSSp:�oG-,,b{{�	�D6����S�N�ԩS�Bx�+7�p~�����Ғ����������x������T*Y]Y���(�[��E�x9���aaaQ��Pȣ\.�T���|>q0��3�����z}�5�0������L���Q��J��w"&��I xy��h$��� `B∰�}tJ ��w � �q""�����Q�T�L��p�x<��V+V�B4�����    IDATM��&����F����z�p.��vۤ�&_6�Q6�OM���r�Ċ&��ޮ�Q��� O �͘X�}lnn*�'��汶�jbU��l6�������}�h����O�����ʈh\��e|�+��+_� 055������/9^��W�/})<��Un�N�VVp�3x���跿��M������K}l����J�{�f������U�����&O@���;��B0 �R)��h�T��s:��D��5lp7��i����Lp'��|l�R���CDd�����82Rlp-�'|�_�qk�!"���)_�
��b�܉�(�J�v�p8�}�r�x�k�J��f�ٷQI�4D�Qd2<44J&��cǖ�>LO6P�RA�RF0�������G�X,�T*!�h������u�:SlFmcc��sʑ��d�d���D���}���p��_�G����/�+�?�𲗽�S��B������<��Μ�w��]�j�T7"��p8���9�v��K�VL���SL�����M��~ff�_��t:��PM���y�E�1h������$�r�{�F	�ʋd�n�S9��n�x��Z�:�N�����]�����^j�?[]��9��� � ����M����p8�/i�B�&Vt��bql1�貺�.J��r\h$e���
�<R���c�8�T.�Q�וi'����5��|���8~����T��
Fhcc�]w}���������1�*{�v�XY����r݉'��=�n��w~"��Z��o}�[�ַ����-��ꫯ�K^�\u�N���_�����6V/]¹��q��y<��8�666��FD'N���i�U�.���j�T���bq�B�T���;��F!���(����x>�!!�(�a�������ɛ�i�hT��.�\'RP�e���.}�'"����� ����`��y� n�O �o �(""�"�B����Ԋł��=�b{{�Ċ&[>/7���2�},,,�}�LNa}��F���������SSS���!�(��{8~�8���͎KKGؤ`�t:�|>��N���p������X,�̙38s���7�˅cǖq�8�|���XXX���"R��p:�V|p�n{��������666����g�y+++�(GD2??�H$�\S�V��Ű�,-���;�vv�M��~���z��B�`R5�!��7��J%���iϵ��NF�D��7 ��
���c��J��ImDD#V� ��Յ���� �
�� �bq-DD�Ajlp'R+
P�%J��4�\.�|
��v��g��}u�{4���A��4����l6����'�����e���躎��\uՉ�k�� ��r9�.��sx�+~@����.�j<�!���m�?�ϟ{�3�ۍ��9,<��}nv�X������aur����2��,���<��<vvw����͍^C�������n�����.\8�i&	H$��7���6����9�!�s����`��)u���>�ۍ�r���|iϖ��
�z�;D��դ�S~�'"�"�x/�o6�ȱ��� �
�] �@��r���%�7�O縭>���N':��ե�%i3������@�Z�F^���X,�t:mbU��Pȣ�j��v�Y�!�H2�`��;��X,�׋F�abU������G��������w���elmma~~���Á��>������Ѥk�ZX[[�ښzZ���D<G,G,�k~w9��p:]p:>��������l��l�Z�RA��A��A�\F���5�����{�L_'"+\u�U���@��4��wd�,.��������0� �I&�������]����˅hTʓɰ��H�XLy~�l6Q�VL�h�y�>��7��X,�V�a���.a�I	�lp'":��������d6�[� ���?�߰�"�C���*�w:��e��M��D��E�G��B�ZE ��,����@�|33�}��bq����:�ٌ�g>55�w��������t�Y�azz���;:�N����m,.�ёH$
�P.�M�̾VV."�J����]�'�JM#��3�2"��ߍ��}���ĊF��wB �v;�p�efq�=���Q����焣��M�JET�U����d2�l��<{9���ŕ��y��IJo�T*��J��p8����.cl麎z�.�!"��<�V g�.��V@���_ �nq-DD��á�3�85iC����H����$}fK�.4<)�*O(�� z�r�����t�2���f��¢I�P���ŋ�u'N\-&���4MÉ'�u���b�gaaA�����Q⨸\n$�����.��G!�T;�f3b�'g�����BA}Adw~����Z��P����_�� �1��������� �c �
 �Љ��J� �DA ����&m*󒈱r9�gv ���ML#e�Yq�3W�����@ �P(dR5�S���i33��z�d���
��G�3� """"X\\�;��*���Lm�Ӊ���B� 2��MOO+�t]��܍�p8ċ��c,�׋@@}>$���p��6������-P����H=DD��q �hZ\=��� �7ѻ��k!":�
lpW
p3�HI�T��L�6P�QGlK�]4�N��\N��455eR5�����l6�k���te66֔�5M��ҒI� �;���������)DDDD��|]�}Gc�Y����v��k��>Z333���l�Vˤj�#�+�Xu]G6�1��ɗH$������,I�s:]
�S��D��L[E:[#""Q������B?����1 7 x7 �VG(�y�^�K k�Z�V�����!��X�����n�LF�d�H$��a0]�����Y��R�$&��������TU*lnn�4�<y4��6������ɓ׊���v��j"�Á�E�%�z��L�)֣����;&Uc/R�B>�G��6�{��Xy��X�hD���l6P��M������9�WE��$�٘� �� ��C<_:�/ ��PG��P���nQ.������i"Y�PT>�F�$k�\.�|����k���z���v���<ҡ���F2���QZ_W��;N,..�T��K+h4�[�`G�1�""""��3;;�x<�\��q���*"�w�Y
#Y__cs����+���md2l�5�&��b��4MC,��;�ͪ�hi8�ު4I���4M���w)���!��.�1���@�LF�bw��� � ?�^kK!"/�������:��Μ.6�I�Ѡlp7V.�W^^r:�����j�XT_䐒�hx�J�rY�fnnΤj�)�ɠ\.)�,,,��r�Tu:\�pN\w��Q�%&""": �ǃ��:!�[YYA���%�h���%�%�f����m�*��Á��Y�tzOܡ�E"ax<��ilp7V4U�u�z�<�Ɣ���N����9eV����TO�f�;�d|���!�k�����x�[�4��Y\�ؐ^h�lp��D2is9�2Q�@�n���s;W�Х���
S�i�*��9!Op��I)�N���&UC �N���$�Ák�� ������q��I�g�X��֦I LOψ�~����dr
n�[�f{�Faj*�|^.�Q��M�����y�P@��1����p8�D�k��"���Z���;��DD?Pp'�� >	�_z	v�>��: 7x��Z��,'7�3i�nR�J���ߊ��7�i8�\������V>�z��(]���ؠ %�ѕI�Өժ�5��Kp:9��L��=�v��\�D0??oREDDDD�_2�D*�n$��.�y�)&<�LJoo�[�t0b��J��RI=��F
U���hxRx��7KÉFcʀ�v�-Ny$�;NrT��j��lp'"B�g \�?���C���W��p���BD4����_�ղ����뺘���M���ٌ�y0���3�{��j�T*�5R#��n����s܀!]ױ��Nqw�ݘ�c#����&VV.���������r�p��׈�����wC2V*�B0T����dP��|>��꽽��-����p8�O�N�ɨ'|�p<B��r��7KÉ�b��B�ˈ~?�U�uu�;��u|�� >�c�)6�n:���R o�Mk�!"2����ss��jU�XJD=�Ei���S�V��É�:i���N�)�OO� `��Ѥ�^�WL֢+���#~�,..)Ӷ�x[[�����N'���Z�*"""":�N��^�W��Z�bmmդ��9KKG��;�677L�ƞfg����v����1� ��V���jU&[L���h4x��`R8N>�7������[]�X���'AD6��?�8�w8om9t�xB;� ��J 7 �{��߉�&^��U>o��ܐ��D���#��N�I��C.���w�I���hĤj�#�ω�Ҩt�2��ccc]����bff֤��9��=-~׏�㘟_0�""""��'��໬�g�yJ��E�J$���5[[�hq
��h��l�{�t�vۤ��ejJ=-poO�WEÓ�T�Y��,��t�����~"��z}H	���OD6�p�� x��[[��&σ ��'��G�]"�x��N���S�X*Z]ѡP.��Y��@$5���'����g?�Z��RQ�b�R�d-:��u�{29��cR5�����f��\s��Q���V�au�������DDDDtn�'O^#����D�P0�"z��G��ϻ�.66��>J�DB�n���eR5��D����k�0��i���i⹜zO���Ŕ{حV�]D�`0`u	c��h����}��l"���O8�} ���2��M����G{��p��&����pS�r�L� �����X,fR5���唩N��(/-�N+��RӼX0;;��1���1=|�z�#R��OL�#㭯��T*)�8�N\{�u�|""""�W_}R�,�l6p�ҊI�s��$"�����m4��*����y��z�&�	���R���^��D�r��>�u�i����
z�\�������R����s���&�9 ��"�ش�6�O�u �Xp�/ ������9V�E*岘TJD?$M���oh8�NŢ:=.W�ԥ�I��=/�@��DF��77���Q�����3��|���g�R^z��&UEDDD4���������O�߃�xG�S>�u��k�cS��dR�f{[=q�Njpgz���b�����y��H�.a��j5�K "2[��כ \�. EK+���ɬ}t|������ �3CD����F�˻=Ϸ��ku	D����
��r�L����I�����W�UQ.��ki���I#��� 'E�X��S�=/���	d�r����K����y�EDDD��xp��Iq����A,055�pX�޾���z�nRE�4;;���u;;<F�h4
�ק\�w�I{��{`,�ۍPH�G��|"5M�����.c�U��w)4���9�6��ߍ^,?�l���t�� n �) �) �C���*���md��ɨv���cu	D�J�RQN=�4�(�O��ͪ?�C�<�I�؇t�85��X��f�h4ԣ���L�ƾ666�n��k�9
��iRE����U�J��Ák����QDDDd{'O^�ۭ\S��q��y�*��;ztY�\�u����T�=i�&^^�d2��:"RxB�ZE�R1�{p���C�5�^,�T���l�VS7�ٝ���4M����w":��|��֓�9��Ն�m�޺ �a ��} |�@D����b#��֦IՌ�n����(�#C��l�J�"6�&�Ѻ4��=������e�$.�J��奎Q�t�X_�R�=��g���t]�SO=%^l��8r�IU����y$���3O?}�'^�-��F(�n2���F��nV�+�L&��ĥIktP��R�{{�>k����ٺ)Nu���bq�s���NjTi�ZʰM���ND�Q�= �
`����m��������A��C f �	�d�g�,��hPR����%��=k{{[l%���w��5/�S��M&�L��>��J��rM*�>����5�����ifg��+Ȧ677�j�S��9
��)�f�V+�tiE\w��1^:#"""[�����⺍�q��FA�ѣǔ+t���5������zBZ��@6�ޓ���F����t:mR5�!�J{�4<� �g�;�$X]�X��@p�% ��q􂙧��� ��Ec��t9u ��Kv��q�߿ ��ј�^Ҫ�*��1
���ODÓRUB��8��#��M$�p8�dj�tZ��JMsst���x�>?�����u:1���vcaaѤ������h��p����r�R�8p8�����1��*VV.�T=���4�Au������Iٓ��G<�����Ű��B*�
�ՊI�؃��@"���!���p<�ؘˋfD26��U�lp'�Ck�g � �� nG/�Y=Ɨl��4��>X� 	�'���5�
��q(E�^�����eJ�ZU�~��Xce�9�z��X�Éx���F���n7�GdkkS���񈣼��mnn��T�/..��d��t<��Yt:�*�׋�'�1�&""""�-/G(R����w�n���f�49����r���ee]�b{{ˤj�Fܥ=)^,W^~�u�&���j5^f"8�|~��k�ZM�����h�l���! /���� �ڐ��4�6�3 ��M �`�;��A^����P)�M�f|�;�����4:Tڼ��t:m�r�4��)��]^�^G���4==cR5���dč��(u�r��9�}q�)�V���x�.����̬	Y+O`qqI\����b�Cz�033#��nmm��
te�N������F��4�"{�Ţ�x��5lp7��w����n�M���@錁� ���rA��Npg�;Yh/lh�G/T�3 ���.:���NW�G� n�޹GD��v�⋮��x��L�h��Z-�g�=�a���2�}��d2ɍ�H����T
G��':8)).�!T'3ҕ��di�<�I��mmm� ��O��g�M.�ۍk��N\W*���zi�ы8;��\��t��n���Y�\�I\[[&Uc?��r��jUݬG�K$��烼[�p�36�ɤ��v��t��4Mc�;�i������̆v2��h5 ��;c�hdip�p��6Mq��L"�BR�x �׫N"����Y�n"��I�؇���t���?"��[�v;�5Lq�^������t���c�D/���O�ɊN��]w=/B�ĺ�k�K��Ng�>�&�,,,���)�lmm25����w�r��)#�p805�R�az��"���W�wc�|>�|���|^}�@Dlp�H���%��������$�9��?�^H27�Plp�Q����7�C�ᝈ6��Z������	Ռ�Z���m�^Od�F��Z��\�wc5��J���d���F���(ԇ-333&Uc/�v{{�Cݙ�1u��������r���<�-�j����g�u�pDL�$""":�z>��	�F��r�ȑ#�5���u�*��X,�`0�\������LN���^O�Q.��}�t6P�Tx��h ���o��IO��ND���g��^P6��ȱ���VA�����?� -�*#�Co����K���q5��̙o��n[]�D�F���	�*�)�]J������Q>��bR ��z$���G{ӕ��.VW/)�h������D/��f��!7�9r��>����8~�*q]:��Ύ�ݎF�ȑ�p���5�h���8j�$�V�����0
��uu�O�3��O�T�}H{���&2J��N
�""�B%�z;�kh���Blp'�=��~����� �ZWM�G��:{4|onl`�)@D��6�{��LG0�4*���sd�������:�i����>
���嚅�E�f�vwwP�T�kR�iD"�*���r�rYX�����M�˅�	�_���3�<mRU���^��m��Z-������I�;;��=:8��-6�J!4�A�K�=W��ib�܉dLo�U���j~�!�!���ػIc��4n��ID6��Z�\ƙ3�����P����o?buD%��)'F�j��%    IDAT�n��a+�|�JEL�`���:��x�53��Q���T>������c���麎�����e9=�F������'��v��\.7���%�4n���v�5�����t<��Y���k�����%�K�Vl�b���hZ�⺮ckK�N7==#���Li��^�pY���D�r��>�u�|�Ċ��`��*�N�F��sM��zOD������0bs<գq��c/��NDJҡ��]�p��.���麎��� G{��j�T*)�H�D4<��ZJ⢃��B�07�G$�N��T��_\\2�{�d�ń�X,��~U�U\�pA\�D���lBEDDDD����4����U��Z(����:���M�Ⱦ'���k2����I���̬���~�/�M�+ez����B��v����$LpW�V���KeDd[�oh ���Xc�;6?��>��a�;�"�ܰ/m�<�M��O�F�c����ޮ�eM�\.�|�&G�I�ՑH�Ǥj�#�͊M��A%��w����\�H$�L���.^�S܏?�V���D:-��--�(""":�"�(��'
y��^}A�Wￓ������uf8����,�n�r��G����.�p���A$Q���s1+%I�s�L��z����%��j��|�w"PE����kdgC;jlp��.�^����� >6��Ұ#�:�|��Q��Q�O?u�y��2�&V6�Q>�#���X,iNG@�u��{�5Ҩi:���-����I��[�TG���H����g�# �������L������.��]w����j�p��Cqb����X*��wm2�&N>�V�l:��Yu(B��B6˟�ђɤ��E��F��7����v��C(�3"|>�N��e��A�>��v� ��^���� �Fwu�јc�;M�= _ �a����w"�������*���~��y�˿|��2�&Z�XR6[k��X,nbE�O�u�`j������z��L��^���T===��&�x��(��|N�Ӥ��Gu:�=��]u�����׿�ň���0�p�u�pAO�ٳO��h�R]�6P����j���)��~��������i�%�=N2i�4���E(��.6��T�l6'��h����%�=��]�%���F����?�^8�WpS�&
O�h������uшt����V������$�s����7'�FNӝ��.�4:7���tJ�"*��˙u"�����������I��[�V��ζr�������*��)�˸pἸ.����kL�������,//�ǰ���$j����"+�d��r9�*�7)���nawwǤj�'��s��7���D<�^�d�{�4�D"�|��v���lpWi��h��1k�������a�z ��N��w����?�% ��Æ��""�� *�
��4�iuR������3�~��2�lC�+mj���,���8�,����܀\ �$��` �*Y��fڔ"�i��lSmʔL�-c�v&��LD;3ӭm^�'�yݣ!�XE �;�{"��;FV� ������!�G�D�y��|�a4�|]�u���$�Oq�D��\`���s�����q��+����f���C 099ea�&�����RPbd$�"DDD��"�����u�|{{��7DWr8����T����V�O�088(�9::�~����C(��8;;S�M��B���ψÐ�k�ui�K�;'��w�RI<���*�����h�t�5"���F�.�O��9 ��x��\[Dt7�@�Zſ�����n��Y�^��������N�B�SZSW����v�����5��)�r�Du�[��$D��;�����ts���םN��+R�դ+�u]�l!�mnnHW����)興���z�^/>|$���jx�n��;lzzn�[X�L&Q��D��I��v�0p||���ޣ�����������^�h�@  ������irs����á!"V�:��Nj�S����q9�^�\kD�ǀ;�e��x�0�gh��:�)�l6�o��G����oh4�nG(�����qp���V�zN�^��������t=��x�n8�
T���XlTQ7�'��H�[��o~ɏ����C�v�*X ah�Ú�&���
7 �˱KK��x<�:#"""�s8X^^���T�x�~M������׏��	a�a���"a���,����wc�H$"����@��t ��l��O�Q����F]Q7Dw�����^ {F��Dw��@�ߢ5��b��� ���&?�Ķ����.��c��c�h���ݝm��?�=��x[���S���۷o�����(��w���ur"^-*;ܦ��f��C:����6�M�
����W�M�M���G8���Uh6���ٖ�-,,��:�X,bccCZ�v����M�1u�/�X�������p*l��_�^����C��M�*LLLJr�Mit;�ؘ����ST*D�n�`Hr��D6ˀ{��΢s9�3"j���Y�T*
_g���k}h��h�����'��8>�#�����)��?�w ĉ"R�4Ͷ��.
����_�o��Q�������޾yݶ0?�L.��>00ha�]G�^��i^X�+ꦷ��i�����'�H�^O{jMq'����C4�� FFFuDWI&8>>��~w)��������g��'��)���\<�iCCA�ϫZ�2P���锞M�rYi@�n�����x��l�����L4�?��6s:��܉��z��n���j5��yM�p'��5����@����Dt	�D�����OL�S��7 x���ڽ�loo����˗�ѱ��x�����'���/
]�'�ugg�����!*�7��i��H�CQ7���lH��GFb\#j�h"?�!P�Q�3���%��������N������S����q���'�)cffFZW,��������i���_����B��T����Iτx��N�W���t:�����t����/
	�B��:ι����O�����J%��|.C�q�������5�[`����>úx�x%����K�a��X�o�����C*���&t�V���&���������l��J���i��U�����]_:-�����B!���DB��x<ҵ�tsGG��)������)R)��a�ۍ��)E�UL����[T�Ui����4"""R����/� 
�@�����[��@,6
��/����C�t��Ok
��y�K�i�t�~:�N���	��&2�fk7�9��I '*����sH�D�̀;Q�����r>��[�ڈ������W���s ��������d�&��q���׋��i��O �@�ow�R� ����� ��G� uV.�C4z��W�ۯ^�#����G���i�t}�|�RI�.4E6�fv��jH����h���(��
;�]����'&&��Q��g�I�Zkko���s��K�4,//��_��)�r����N�챝�w�V��~N�����*k���=b�<����p_Q7�)
K�x\Q7�Et>���j5��o��`P|���qh�~?�������v�#"l�=�?�� �:�Q�`��H���w�# �>��9&��MT��K�޿������t"�"
!b`` ���+t�@�RF�XD>�G���l�|^I�D��Cj���χb����ސN���p8����v6H$☛����p8��Çf69<<�5M���66�vջ��
�1==se���x�`o�|��1�Aggg��X�_<�9�.��<��W/9Y����l�i:��V���/������.1;;��-�I$�8??S�Qo��]X�Z�"��0;ɦ���%����G���x�8������-z0��qc�>�x#N�3MSz�����b��� 8�l;D��w��1 �~�?�� ����z�1���uGtǙ�	MӔ�Vn4H$�H$.O q8p:�p�\ Z_0���:oS��Z�bAx 
�po�L&��\����Ba��\�n�d��sW�ݷ�Qǰ������P,����!b���vQ��
��{�M
컲&
!�pxH&��蘰���biio޼�gv"""��Ç_`hH�( ��`o�߳�A �~�l6����V�E���K"GG�0M����v��!kNo�G8����u�4��0��n�����������n��6��*��0���:�D���V�� �	 W?u��w2�jM /��O D |� ~�s��M��os�f�j�B�B�R	�Z�A�{$��	_�v����u���	8�ռt3�Z٬8��z���x���񹚦阘�T����mypeaaQ��������ٙ�+v0����������WMMMcddDZ�q�$����Ӱ�p���������L���i��F����nzS,6*�wa�&�Ʉz��4�ϣVcк�dg��ͯD��r�$�H6@K����~P�,��� ��S��2�N�E�#�GD?���_� �$""���������Ł�G6�]6��nN6q�����B��|����p���\.>P%�JJ��G� 5��۷oP������W���H$���Yi]�Q�۷��h4tE2ccc�T*e(�"�(|>�������l��
_�f3Y���Kn�l?��-}/��!�����e�!��-.�g����� �J#�b������ ��)��{ �'�D=�҉H���S�C2M�8���tZ�ZZ����t3�\�JEX3:*~�I�#���LLL(� `cc]��srr^�WQG$R�����[4�Mi����B!]Q����#�6_����շ(�y��\.ff���6aW�WP{MMM	_o6�8::T�Mo
���_X#�@7��>L�D&#��H�����:��9���
��w�RIpg&��]���r�}�sm�u1�Ntw]��� .�ŉ#���D��i�҉,�HDQ7���h��$/���襛����F��\`�l6�B�\X3>>�ө�#*�8>>�h���Ň�:"�b����U�C MӰ��RDDD�}}�XYy]�o���D>/��K���/H��f2d��M�>�`��x�r<~�z�����$rP�Vqr�i�v��}��'��99��"����l6��)�E��5T��+_�4����>�Wp9о�����p'�?>�� ���W�%��t�ouD�F6��
�,=��둭���p8�C<~,|P�i:��Gv�{dS�'���uC ����ZM��kpp��6�H.��Ύ�|��p������S��W.��?���� ?V�Y188������0���aSQG �����������nz����H$���@��mc��S�>]w �pj>�5��gm���mD�\�@�/�{1о�����͘�#��� � ީ��K����`�WOIh|v�2����]G8V�Q�hM�:֌��)�7��i��%a��ĤpU5�W�����u�����E�-���n7?~
���)�����t]���cx�^im.�����s%��i�u{{{�T�\W���A�C��D\z	�ngd$&�a"��+맗D"aᙏi�Z�@6��0n, �����Y�D�Ȁ;�wR�hE+��K����6%�=ŀ;Q�(�����k���OGDDt�fC�6\6͈���hHCֲU�ts��8���088����c�&���S�].b1�pj�T*�|^�{��vcffVQGd����� ^�+++�EDDDפ�ѣ%ȿ�JE�{��i�]d||~�_XS*�8)\1��v�4�����d�NNNx��&�3ϓ���uE������	�ͦ�n��6������,���t����!�_���v��ħqD���V���p9��7 ��'t/��S}���M6's��R)��P(�I�6�d�����$���uӛ�Ʉ�A���4�_�U��ؐ~�p"5L����*�岴vpp_|� �Ӊ��Ț��D"Qi]�VÛ7��h4tEV���Y�����!�0G����
�7��RI�m644$'���n��)�7�N��L��4M���g�iE��}>��a�3M���3��ʰ]��Z6ډz�p�GE|���`���	�4&%"e�Yq���r#P�M��f3� ��떂t}�i �Hk��a��E��4qx(���x��uD P.��?@���C^>�"�z�_�ZM��,���������讛��������0�X]}�@n�YXX����X��D�5==#�0�������&jP�ץ�t3�hT�Y�4M�0����A�\.A��l6����L�4x��N���*���ٗ�i��]V��@�>e�^��a"��;]�⇉���0Aw�萏�����*��υ5��t}�F''9a��ýv�Ǐ��k����QE���x�Xȝ���g"������$�χ��)E��J��o`�u�����T��U###����֙����U���)芬�!O�m6��ტ� ���t�A:�A�TR�Qor�=ҟC"�]����_?9ɡ���v��g�ggg�.�Q�\���b�bA�:��莹�A��A#"��nGDV�����D�$n�TJ�rwhh}}}���-�r�������87���0
k<�>�b�h��a4��Ö�njj^�x�;�uvv���UK���x�����~P8�Ç� ȿmmm"����n�r�0?� ����A�VU�}433+�98��v����I�zL��"��x<	kdg�t3��5��Od���t]����+��@� �&Y;��9.�c ���܅D]����H�L&-|����km��d�l����'�����n���;lvtt�F�!��w�2���᦮�X\|+�'R'��bss�R�����%�x�h��E߽�])芮ca�\.������?;��S�s��t�"ݎ�m}�l�JYQG��������f�)=����������Ȇ��'~���-t=�wf �˔�ʐ�5ZAvډ�-�d���%�`���W`�J�b���l�)]�a���b1E��+-���uӛ���5n��?���\�^>��ؘ��Ȫx���:M����#�B!]Q����x��	��6�JbwwGAWt�PXzI�4Mll�3X�����{{��7���a��a�lݜ����A t}����r�Ӗ�,�4�-%��:�U� f ��J ��V&�b����
��:��+��]R�x� ީ8���T�Mj����$�	����^���5��CCC��8��N���h4�C0���-m�}j���?H������������ h����*芈���U?�<y
��)���O���{]�u8<x�(�;8�G��)�*"_*�f38;;S�Q�_�/����Nu�[� |>q(��wX�>��N�'�����ٽ�lz;�����~��O�ʄ���F����TI���@+�>�V��W �:��+뀉��Ep���V�M�89�K'Z���'�����0�t(N��W�����x�������Ǐ�ϋ�;N,.>T�]���:NN��]w`e�1'P�(�ǃ'O�Y��_(���۷0MN]�6��s���֔�eN	� k���t���~��b���8��##���ZUz�@���x�5���� }����=Qk[���@���QG1�ND��@+��s ˸x��`_DDD�vzz�z]4EY�N|��0�J%���#<��I��@*���b1K��掎Q��7?NNNq�{lllH�ƆBaD�Ê:"��������'A�\.<y�T�"""�������� �r	�_�F��P�]�������������^CCA�5�t��gv����	���D"�	�v�4Mzf�L&a��\�n���z���D���sӫL� �����d���h/�h�t�5"�e�Q���S�}�8>�w:��|�@D*���\.+�a���h.���x�5���ѡ�u]wH'M��4�MKS�e����咥)�,��▏_t�h    IDATn�l6���k�J��I@k�۳g�r'""�N��?����V�U�~���R*���:>|$��[��C�533#�0��������t:1<,X7��tS�`H�%$�����D�g�����Y�i�J��J�,�!�����?��@��?B""Ep'�nu�O��9\�s�$]�i���KDJ�V��ANP�A�T�N�`��>�Bgg�V����v:::D�&�999�i�pp��B�\X�r����PQGt�z�~�-*����O�<���Q�u���ē'O���z�_c��7;;'��P�հ��AQG�Q(�����&�JKσ��FGǠ���̣�#E��ٙf�XD����t:14$��͊��'>��Ψ�H�XNh���P��|
�� W�QW���3hMy�Z���εEw	���J''9�]�9I�&ɤx�{8a��F������k��vÐNqw:�����ib}��t�l$��Ȉ���:j�*^����|�j?�={&��GDDDw������c���6�oQ*�tF�588h������������Y��ibo����allLXqz�g��&��HXX�H�u�[B�04����f��=����_�uŢx�$���E���0����iUDD]�I?"�������4Z����; �4�V��Q�J_��d2)�n�Fv�[��4�9>>����u||�jU<�}bb��=:�P(��P��eaa�w�r��ׯ��n���������3������Ti 0M��oq~.��C��p8���#iP(�N#�I+�>
��_"I�R�<�@8B__�������F%��M��)e���9�l�]���;�B��V��&�5����@�@�_�5L4߹ֈ�n�w"�/�����S S�x��tR&Q�e����p�x�/]_�^��INX#[�K7g���caM(F���(ݎa����8�NLMM+�.���E�\�8�N,.>T�]W�Xě7ߢ�lJk�^/�<y
�˥�3"""����x��1�����M�{�&��J�377/�~�h4�����#�D��̜��4M���i�Ǎ����j5^��l���ɉt�]���@($����duCt�i�����6��i�(���y��.����	�a �h�~��E��^`�����	|
��@��}Q���]D�T&��L����$�I�냃C���S�M�9>>���i&&&vԛ��8*���f||�-�fM��Nz3
ctT��:���kko-=T���x��)�&�q��cy�1����M���G:��g�
��o��ܐn*����F�S^����+���
��5��G2d��#�T�L&u�[��t��H�i��f�ؙ�*��'�7E@�\�5j�����v1���oUѽ�OD�+�A� �_��H�z��|^��M��n&�I��hk��œ���j��tzQ,�4c���|���똙�Q�]rvv���i���7t�\.���U��<�r'""��t]��Ҋ4�����:�]��t���/�u�L���=�_�ꬰ�4M�퉿�R{LLL	_7M�D\Q7�������M�f�S�m�_?9ɡѨ+������n��
���:���9�(8ؓ�z����W}�Ap\�CDD6H�S����0��nz�aҵȭ�Cd���C����dj�8*���fd$���a;awwŢx����Ç� z�M���f���fiz��� �>}�>DDDw��;���ᰵ-l��{v����mV�z���:���l�Ǐ��w���n7���!�t:�j�����32"ґɤ�l6u�;��R[*%>�'����N���dg�t�}�1��$.�y���z�DD�`W�ţw�N��."R-�I������t=ɤx����ࠢnz��iggg��	N��i�����h����yE�E�a��{y0zpp��㊺���d�x�n����ߏgϞ��v+茈��n��h�ۃAk�۷�?������6�ሥK��j
:���N'���Û�&��v�4�㬜�ɷ�����%�{D"Q���i �e֐�*]w���v���W,�'�3�p�l�;��IS�h�5 �)"��$��5q9���_�x?�\kt[�at�"�1�z''�� �)Ht3�|^:=*�q;�pZ�F��J%q~~.�	��
*�.*
��ߓ�����!P�K��X_@������ɓg�u9�ÉǏ�"��Yy{��m�n��rcq�.�L �o�#{LO���o<:<<���l߳2��nnttT�z�VE>�9]v�F���s����n��>��M�J�J�"���i�w��@�Z�����M�A"���;�\�K �D+�F+��� ~�'ww'��j�xUi(���T�M/1�����p:�wo�t:�J�"���Oe����ޒ����)�~��ޮ���;����ϲ].�Lb}�=���}>�={��ccDDDtmN�O�<���kww���;��Ç�K��Z[[��:��<���۫��:��Q!���_6���>�Ѩx0D2��4_8�N��^�"��@ ���^� >��;)��͟���@�|�1�NDt���p9��{ �εFV����ɤa�WOU�u�pXaG�#�_�u��Gu�{L��ёx����C($~`D����qr����Td�4���;��χ�Y^D�v�D�j���x��9<�>��"""��p�\x��,����boo�ަ����'G�u�����!��s�K�{{�h6�󱟆��IaE�\F6�U�O�����$�O��H$"�]d�ٌ��@����^V(��3�p'\��Ck�� �v�-"���w"��k�S��� p9�.[J�q���h4prr"��M㡛�T�������x�/�N<~,��R{lo�l�����;�T*Z
EMLL"⥨n�cccV&�����ٳ���뷿1"""�r��x���~kS&��v���csWt[>�ss�Һ��#�r�v����ȈxA�R��񱢎z[$A��;����|硛�Y���Q*�u�[dg��\������t����ddwf�R��+�h�D"�6`�����>���{W�M�$"�C:��
��t:u�[dS�����]_�ٔN�
C����:�]�B���wQ���c�:������LZ����5��y��1޽{g��S__�?�߅DDD��ׇgϞ��������p���:=Z�N�T��]�Nh]@_���� ܒH�#F�hԑL&u�{|>�tڱ�̓n��t"
kdg�DtY ��/2�J�F���5Mcơ;$�
����(>�W;�ѽŀ;��>�� ����εֻd3���-���t]��&��/�I�^��`�OD��9<<�<9�]���m�A��̌t6��4M�{��fS<��v�/)�n#�J�ݻ5K!�ִ��T�}����ٳ���Z���ٶ���:onn>�OX��,��fSQWt���B��������RE���{������H6|��h �N+ꦷD"Qh����@6�MD����\�p.|�ن�I��D+DDD6�; �ze ������5Z��Z�Z��&�CD�n�F'''h4����bR���fxx��@�]�ժ�!���<���zWk������r��AU*elnnJ�B�0���tD��N�,�ܝN'�<y*�Q{<{���w�����gsW��P��Һ��]���*舾O�����j{{[A/ ��S��Ð�-��麎��aM*��a�����a��\V:���.c�]�P(t�jI�Z�*���@������ڊw"��+�l�+0𮌕p	Q����PN�SQ7�%?��t:y��f��5McXW���]4�qSS��x�uD�K&ҋ9 0?� �ϯ�#��t:���7�V	�++��Չ���=������3�\.K�[[�8<����r���|����)/,tP,��/��rY�����}}}�D�gd�T�]�%����'��:�f�N'��!a7I]�������6��,��l�m����|�� �3��U2�ND�p'"�>E�p��o �@�c��#V�%DD�ɤ��4MG8Q�Q�(�8;;֌��*�7
������18��o�F����}a��똝�S�����T*a���x�h�+j�l6��շ���hZ�g+[KODDD�G���S8V.��X_���C����x�����@U�����ֶ�P�9�=M��pz�*������c/����9'��$�BӮ>c1�&�٬��>No��T*h4�f���@�>eqh'"�B|JD��>�����r��% ~��!��H�f��\.'��V�$q�냃C�z}���M���P���b�S���T�Ua���uD�����|���W��V.��۷o�l�W�k���Ň���V�Q��F���b��4M�{�N�������$�ᰴ���R�����B"�d�W+�2�\�bQQG����CCAaߋ�#;��fs����'��
��יi��āvfm�������~o�"";�V��B!�
Z��T*)} ��uӛ��,J���frr��
����i��܂�n�*�����ߓ֍�O`xxDAG�''9|��7�׭-皝��Ç_��Q��OX~5kk�H��
:�v07'�H�L&�s��~��Ok���]NoWebbB�YO6��nG6��0�޲���^.����e����g�]Fv��g��rqx���DDwSDDw�(���Q'd��*AM��Dv�;��&R)�C�Xl��j���X��n���
�D����0ap����vqvv*�[\|�׫�#j���3|��+�&��b�Q,-�@��a"""�4,baၥ�f���o_#�I���������24M�ݾR)cssSQW�C���g0����?3��8���k��"NNNu�{4M��H�Rh4�:�-�HT"5�&r����>��'�8E�;3B��VF�b�� �M!"�������y�}������L����l��ūP���c��.���
s��d2�Z�&�����T%L|� t����AD���w���l�`;,--��R*��7_�\.[��D"x��\.�͝�O��ˏ�Ώ�����k�9���OX����N���34�x�V��K��>cc�p��[%8��N�pn�GX#;ۤ��m��f���Dt���@�[�z�J��8��L�%%�p�������>ѝç�DD�_�o�)�� � "����2��x�3�f��Τ�0b�1E��&�0�����y�C���S���i����S�:�R�T���!������_P��K�R�7�|-}o�(��/8������n7�>}n�Bs�=����h���S���YݒD��4��-��[�*��:&&&�5�j�TRQG�Iv&Y*�pz��]v�x�044(��������
���2���hsd������;!QJ���@+�>�V��W �:�WGp:,uB6��a��i҉1ts�D\�z(�N{��9>>B�.�J255���*|��)���
���Eg%�I$	i���8FF�r��j5|��+�A���~<�����DDD���ߏg�^ X�/�J�曯Q*�l��i`` ��sҺ|>���=�Ub�Q�|~a���)R)�IU��F������a�==/�V��PHX#;Ӥ�k��\}�l6����5Dt8�Nh�@v�����4^��)Z��ڹֈ��p'"�$Z���XF��y KD��l6��d�5##1E���d2)Y�at�S���l6q||$��z��&���־
kt]��켢��*��떦�>x���F��7o�E.g큹��'O�{���Hbpp/^|���~K���g�曯Q�27q�8�.<z�, �j5�{��3�r8�����T����R���s��m�Z��j����	���a��;݌l�L&��� ��8�������y�=�֐Ə��J�Z#"�n��;}.�ˁ�1|
��t�/[��DD�I&�+}}>�~�4+��F��L&-���G�JW�OOϨi�����ZM������������U��Á���CQg��fo߾F<~l�^�X^~l! DDDԛ������S8�.K�''9|��7�mS�m4<z�da㔉���P�ՔtE?lffn�[X�H$q~~��#���98��i����QaM&�A���_v��|d�����w�r��F�q�뚦���ߋ��?�DD$�����)�>`�ﻝk�}`$�N89�I�r��}�q��)�˅htXQ7��ѨK����~�zfj�f����mi���D+��~�r	�u>�
:�v2M����`��LO��ѣ%~�!""�`ff�-[~L$�x���"!u���iK�wvvprr��#�J����f���럅�4LL���7u˗p�f��a��a'��Gv_�U���uCt�N��������eۉ�&.�#�h�- �j$""!>�""��:Ƨ��,�y ?C+����n�|9$�;�4M�R�)���#�e�|��bQX311����uxx �@�)��$�	锼@  �*F�K�R���c��������;�k���G���3�\�i�DDD�������ʵ�G���b}����]��`���:��a�N]�+�4���v1N�V%�J'W[��G�#��Q.����4M�9I&���@tM��^�\ֶ(��{p�h�[��&~h?�\kDDt1�NDD����hާq9�~���,��u�l������PPQ7�G��\�i�Z�&�@500���!E��֖�fnn�(����&
������E�.����޼���ի�/ċ/�""���������D���M����k��ݱ�3�C__=Z�j�����p'E����J����;�H�ޘ�Ooo68::T�Mo���ִ6 �w�B��n�Eq�>}�� �"eL�D�(>۽#�&�5��!?E+��hM�
""�܉���.ާ�
�����ʓP�0��h"��
��t��lE*�\"��e������a��)�SSӊ����S�v	�Ӆ��yE�U����[��1]ױ�����w���	^���j�R}__?�?��p��Έ������ǋ_"X�o6�x���I�g_�N��ciiEz��4M���r"x�9��/H붷��[ި}B���w���kn�f���$��D�k���ޭ����q؆\�X~��4�[?�h��V�7 �r���ڊw""��6Z_p~
`����`_�0�ND�"� �D�p8u�[�ͦ4��3j�j��T*%�	�B��*t{��`���بt�ٯ\.c}}]Z��x���M�1�]T,��7_�T��P��p`yy�6wFDD���G�����x<���*^�z�\.gsgd�֖"�wĝ�m��rhd����J�}��y��iE &`�����tbxxXX�L&�h�u�[��r8��]��;�]Ђ��s���U��?h�*""�UW�#QO��(�ˁ�l��b���:%�J
�:�����d�t]��訢nz���d��9�]�j����}i���C~���t�u�b������S�١R���_"����I�4��/�ѣ%�:/����i���{�����P(�ի���z���O �O�f�88��!{�|>�j�4�����#���!�/�����~`���1����#��}��h4*��`��t�!}_ �����8��a]�� "��Ā;u��/H\����Ư(\JDd�j�*�&622����S*��ϋ7&����@�f�RI:�-�r��B���(�J��χ��qE����&NOO�u����뷩{5�M����VP�5�����m쌈�H=�˅Ǐ�brr��I��x��kT�U;#;b~~^ZW�T���NAG$���(=S9<<@�XP������u�4qxx����5::&|��4�6��������_�0�ҳw�0u�S^�g &p9��Q���p'"�n����|�%N ނa/Q��V��A˫���d��<�>��#)    IDAT��aE����w��iNqW�4lmmH�fg�������������a�"(��`�&��?`cc��%]�ߏ/���`�������x��+�A���`kk�0�������n7��V�i�G��a`u�-������*��(����5�j{{�j" ��PP�sI&�T*�:�M�p���Ȝ�n��CC�-�3{"�a�[����z���=��b�}
���7""�*�Q7kX��X_�Z�w���k��ʘ�����4�M�Cv�Ü�n�l6#}h�)��+
����-��'�(trr�t:%�q8���OP$��j5����4��}t]���
\.������1�����-�ӅǏ�\k�-Q7�����R�ax�~�� p��]��:VV��vKk76�Q(�+�D�N'���u>lJ�Ĩ�fff������}�[��f��&���j5d2�m�ts���W�j6��f9������y�hA�p&|݆��6��C+�>�ˁv�l!"���$�%M /���{���_���εFDtsV�e+S��L�D<~,�	C�z��:�]V����hS{mmm��hk��G�5=��svv�>H�������27�q��y�z�R���#M�077����p8�6wGDD�^��=Z��;,��z��ׯ�E2���;�ۃ�䗝8q�K�����_H89�!�f�W�P(��A���t:�r��w����~�B�s���#����4�0�LF6���~��[s~n�e�8Z�`�@�O�*�[lDDt�0�NDDw����� �3|?�.����O�$"��������W�M�Ǐ����n���3d��)�V�R��j5K<x�m8]����D\Z1?���#�S�\ƫW/qrrb�τ��x�^���Έ�������ٳ���DR(������� ���'��J�����&�S����f�a`kkSQG��lh�i��� �vZg�W_87M���z��@` >���0/K��r�z]�Q������9 ch����wIDD�=������.���x�= �E�49Œ�:����ZMX�)�����ҵ���('�*���#���Ӧ�:::D�X����cbbRQG$�����s�]���	^޹�޼��0y�>|��W��Q��A�x�յ�2�T�^}�j�jcg�B(�t)�Z�`mm�ӎ���ix��!D�] 88ط����#c`@�	!�J��b3]w ���)���hdD<��Z�"��9��r:�܂k�lz���V>�&�)о�ˁv�""�;�w""��.�  I���G��SL�D*%^�><<86:::��p8�@��
�sd2a��PCC�U��>�ibssCZ7==���~��aX]]E�^��.,<@0�Ow�i�������U�k�u]�����G�u��]��i���œ'O�v�-�����ޭ�0��R��z�x�hYzr�Ͼd���	aM�\��>���6==#|�5��?������t	k���g�ts��!֤RI^�"����>��@6�䊿�$.�G�)о������S|DD�K>�� ����AD%[}�v��u�{��NQ(��gpұ��� ��ff�k���NOO�H�G���_(�d�N��4KK���焥� �N�ի�Q.�-�������+�v"""U\.7?~�]�ZH�^�_{�	u/�˅��'p:�[Ԭn/"����Y�����&�P�}�D���'�	�˜�n7��b�P��驢nzO(�^�������ƥ^&����Yn
�@�/���@;�,܉�������f��lKD��
��Ţ�&U�Mo�Mq��|�d�@�XD:���g�����t*���Ou�|����uN�++�-�����|��f��0.�z�x��KsS	u������O��a�P8��_�NNNl�T�4��+��C!��+芬x��!�f�L&�l6��#�����]%���`0��/�9>>T�Mo�YY9�'���4M����R��F�!�1�G bh����>�� "��ŀ;�'% �����CD#��D,�g��K��� ��Ĥ�nz��Ύt���윢nhM���ݑ���/���(般8<<@<~,��z�XYyM�Q�}�l6�����{�������GKx�`�����H-M�033�'O�]�;o"ǫW_�R�������I�NO����R�Y12C($��nM|����j��4T�����3�F��T*�����v�
��5��Nt3>�g�Ȧ�뺞Dk8�DDD���*""�����zW2��z5M��HLaG��0���P(�ϧ���U.��N�����S�^���8;�;�N,,,(ꈬ���@>���aqqQAG��i�������[�t�������_IC0DDD���ׇgϞczz��Y�3�a`cc���a���*��S��U*e����i�g�\.7����wvv�VN�0�������vz��듆��8�ͦ��zO,6*��a�&R�����N�p'���u]���V����܉��>�i������w�j5�r�UͲU�t;GG�������|���̬�n�����{i�$F$Q�ɘ�����(����Xl��
�"U2�4^��w�C���^�?���S ����n"Ɨ_�ɵB1�J�~��Җ�;B���-]�fo߾�n_#u��r	k
���uDK�4sz�
���D�4qtt��������3�j���n�����&J�����p���!""�3p'""�L�^���i\�ED��'���{-�릛�V�H������nE��r��dR<9��0H�X�X���|�ۃ�tr5m����X]}�fS>�{~~�PHAW��� �uBE��cnnO�<���;""�E������|�ό�L�������~,--K'�����շ(�� R'
cxxXXc�&���I/�S{i�|z�apz�
.���#L&�JE~)�n&���_X�H���M��n���u���W(�˶77���?(l����N`����������ӥDD6�岨ժ�Nq����ឮ�p��ޞ�)�s� ���ޞt���4���)�X[[����4KK+���:#����&VWߢѐ_t�(⫯��0/Q{���?����?c�&��?`u�͵�Ǩ�y<��<����nmm���DAWd�ǋ*2�(

:��FFb�z���#T��3H����q�8�qxx������?sT�U�����[#���p8��6 �gp'""����K�{ ��e�&���&�dd�����4/��� �n�R� ��;��|�)� �4������}llCCA5M�%�\���u��?��{(�I�ի�(���\.VVca�4�ADDt��ӄ�?!��zQ�R��W_s��=�p8���x<�m1GG�8>>R�Y577/�ٕ�%���i��]�133#�i6������;066.�9=�s3��\.�t�c"�	��ak��ſ�5M�'E��)|"EDD�L���:���x��ਮ��նt;��IN���jE���`��fff��*�����X��yqq���.sxx`)�v����S8�.]�J�R	_�Rz��s�����?����M��}��z������^k�R&��˗�.��ݣi:��W�����''9|����+�j`` cc�-����~���xė����P��uԻb�\.�w����;��lo׃����yrM.�mw{�i�o:����R.PP���"AQt�%�$��Q�$!r�E�pq���o��S��n��]�\�.��g��]k��Ze���m��~%���Z�w�����&ϥ���I����_�ͻ~�o��+���dQ:DDD�
O����~��(��(���ID3���Q��M�|�;�\�r�n�k��,ݨ8�ng0�m���p �6��E�����:s�ˍ��k��}�x<��m�ۍW�^�I�	Ҵ�M���P���?w]��i�DD4�d2�_��W��&o��4?co�=E�bv4+�̷=u�]���q��""��7?�岨���9�~ɲKKˆ1��n�tz���^���ˊE��'�%�j�~ߢl������	�5늢�,J����Q�)��(��:"�o��qA�����(����^��t:�����qv����,--sҴ�TU�����Lf��|]ױ���^�g����z���2���Q�7��i��ůŊ�!"���t:���7X_߀$M�m����������=^��kmD�F���a�������c3���Eя---A�eØ��s�F�7���D�Q��nØ���l����o�<��<�g�£�l����E�=:,p'""��:"�o���aS"��(��T(�MWG..f,�f��CӕͲ,cy�xJݿJ��R�h#���9���Q�vv��h-},����5��Yx��{|�x]�&�9�ǃo��%VW� |џ���կ~�`�|B����9����E�ݞRf4k�d
�̒i��i��}?QC&Y���O�����	3p���xb�h4����������E�X,X��|J$�7��F#T*��Ot� �hCӼ�4��� Ϣt����<��(��Gg��fz��'n4	�nF�4���S|� �~>ȵ����i!n:����(#����iC������5	����>vwwL7$ W=l�y�td����ߣߟ��Ld2K���oM'y���p8���[lnn��^u4���}���_����D�����:��l6��MNElllB�7;��%\^�-ʊ~�ٳU������PU6L���C 0��f�݋��H����ØB!M��ɛ��������:���� �h4��DDD�������h��(��Y'AD�ͬ�Z�$�b���n�٬�A>���*�|95�+++��Cb4�ӧ��qKKK\]� �Z-�C��{;�����,Ȋf��l������|>?~��_cuu�����T2�¯�����\�V�w�}�j�T�2�ߏ�헦�� ���GH?@��kp��E��ސ���E<7���{���e4��6h��\.kQ6�ia!nZ|[(��@t[fM<tŬaS�/ �'��1�6�$��:"�o�n��X"��(��4Q,c��\.N�B>�3]Q�����,ʈ��T�U�(EN�yh*�KM)`kk���
��qQUGG���g���Ǯ���򗿂�σN"�y�v{�����ƍ�8j����#��|��p0�i�\.^�z=�}���������H�Ӧq�>c0��yVW� 7����@�9�zڜN'�Q���R�h������y�QG�۵(����i6�f!�Ċ<���+�(E�RӴ�:�<������לN'./�7*@�����_r���z�yq/݇�ph��@���D�dܘ@��^�#�LNo��l�e����nAE�)��  ��V��@���v;(
p�\��:�f�#�L��p�^�O������Ʀ��p:o���l6����Z�ׄO����۷���p�Ɩ�%M�tIV�$	�_���f3��T*89�dQV�c�`Ϟ�ƴZMN׷���i����!F#�OO���1}O��~F�Ӷ(#����vca�xk�~�b�0�f��eUU/-J������w"""���sA����f�\.AU�Nq��n�kZ��H$!˲Eͷr�d�� #
Y�]����4.�N#���!��������"��mAV4K��{{���߃�ܬ�.�L�7����DD��x�^������as�O麎/_N����C�ǩ�O��fÛ7���t��6u `c�C����tk�h4��ѡE�O��>7�999� �e�d�0�Z���z��~���\.[���í}�1;�E�3yEDDd��DDD&$IڛuD4�TUE�T2���7**��;??7|]�$�ӋeC��^����W,pyivH(`cc���rч�MS�I�=~�r	�}��7��k�;���+lm���n>����6Y�����򗿂���϶�-���������1$Iƛ7�5Dv�]��idF7
�ME����۝fdaa>���q�RA�^�(���N/�>븸8�(��$��d�R�MS-ʈ��1��HW�ͦ��(~gQ*DDD�+`�����o�N��(���n���F-�f>��5���ӕ���~4uT���׋�N��������N'��̧̑�t]��ޞ�g 8�y��v��Ѭ�������͊���2�%�����H$�_��7_{'�,�u��g���~�N�3���E�_���	b8���wP��ud=Y����iW*�P.f��++�&Q:NO9��
���t:���l0M�X6��0��Y;�g��M7����*�m� �}��!""z�X�NDDdBQ��;���Z��i�a*����f6aI�mH��eCWS܍'?>{���3p����i\2�B8� #�)UU������o�r����H�lAf�����oV�!IVW���_��묉��ۍ�o���W��p�lG����~�[��|��s:�<�ۯ&��(
޿�~�������ź�{~4���c�2��J�ҦE��Bq��e��d2eZX}~���ӖN?��t�h�[eC��pz�dZ����*A��h��,L����Q�)?���(��Y'ADT(O�	7^O7S*�L�3,��H��F�h��t�L�g�t\^^N4�occ�l| L�1����������Û7o ��b1/��vv����F�э~�����o���-�""�Q�������n�����˗S��w�eٜY_�@$b�Īivw߳����F�XX����n��e��+�1������5	�9Q���1�(���`��^�i3u.��(��)d��$�͆��(��E�	V]M@��:�����4M5�I�Re3�t]7��d�ۑH$-ʈ>>1}_,/��n�[�����iq�����/,ʈn���ag�E1�����ކ dFE�\�w���D-?�'��_���$ ��=$�h���`yy����z�}�G8=�̩�sfm��D�ú�c�F݂���v;��7M�
�./�dD?ge�i�h6{1�V.��D"i��������lȅ��(�8ϊ�d���3�4�fӸ�W��ӢT���5��"""��$Ig����Y�AD�M�48�N�|㧴{<�r9hK���� �LB��1^��l�¬旪��e����L�(B�m�T.-̌��ϭ^�k:��������X���h4D����Bܴx��v��r���y��*��2��� dy�w�OI��H$�h4�n��"�s��������ʍ>�@Q��|���1�f�=��[Yy����	"u�0���~	��k3����ϟf��vccc���LQ����wdA���m�p0���t]�0��"�2677!��
�<��� #�w3�n�t��f�wTU�Y�ѣ�	�DDD�F߉�؛uDD��qѴ(�H$e3�4M��Ņa���h�7ݏ��/�4�d�􀞦�R��P(�ƽx���eAFt�z��{�/,ı��	N�?�J�}�G�f/ ܬp����o�ūWo�t:�� �%�2VW��_��p��?�� z�2�%,/�L���'N�}�2���>��'��Dӱ��ܴ�x�g%t?��3..��l0e�d
�h<�1��Y����f�£�l6_E�>>Y�ѣ�w""�	����Y�@D�n��h4cR�4XT8]�\���!���:���(
NOOM�<�nE:�3>}:6��,I���M�iv*�K`���x<�����'E��(�����{t:��|$���XYyI��I"�i��"���2�%é�?���co�=vww0��%=d�����M{z��SΈn����ٳg�q���ժ��	�#�M�~�k�Y!�Y2|]QF�CK讄���ǫ�뷺G%�+�,s�̄���DQ�-J������)ф$I4M�7f������ƾn���j5��q�Ĵ�Q��Xb������v-�l~��-D�1����1N��n����4�N�!�    IDAT�	����Б�N���h�H�|�����fc�˜����F��&A@0D"����h�Y�@D4�P/_�F"�0�x�S��#��b�NgJ�C�N/�����rY��pP�C%I޼ykxO �^o��Nt�A�˗�LO>��"�X���a���j��EͧH$jZ�~r�	�.�D��g�ƃ7�75�l�����E)=j,p'""���i;� �p/�X��E"��,�ccdY���)�t�H�҆{.��<W�Z��3/�����r<���~�����o�h���O|��i�Z? �����e����U��D�P�������J��H$�H$�^���"�{��x������U�"ɟS�װ���b����9�H$��>�ƞR��>L9#��/��ct]�����fhq1c�ܣ^�����2���������8<܇�if5�?��5���p��#~�E2����u^�^G�9~�� #EQ���)=j,p'""��.��i���J"�)�eٰ���v�T*BQ��/���f�!�����h�Z��o�~�����=6F�eh�j�&���^�#��R	��(
< ~����D�Uc�(���9�n^���r��F�����fŔ��D�@�N��pJ�=m�kkϱ��ax�<�p8���>}���h4��H$�����$s@*�K�`3�C�ư��fwz��Rɂ���Ȳ��/!I��u]���.F#^/[!� �Y2��f/P�\Z��|r�\x��9�����Ϲ-��DQ��b��pf
�<����eY��4��0%""�G��DDD7 �rFU�e�yu�]����q��u:�Ӌ���ˉB!oaV��j"�L�N�~?
�TU�03�����a��Y��r�P.�x�!�V������̋�����F�����P�C�4��~�-(?��r!�L��t��n�s��hB�,ce�������o\���:r�,��w�j5��%=��67�&�;�ժ�������p���7�E���u<�����s�-Z�|�Ϡ,����s�4cM�pp����)[Yy�� ]�qxx����!�B�Y���i����s�k_Q�{M����i=j,p'""�UUw �W�΃�HUUx<x<��1��l��S��*�aq���D�^�`��VP��T��[�(�n����fa4AQD"�Kq<��>:��E��mT�����>��`0�C�ͯ뿁B� Y���y1���k� ���!�N�f���lr��� "�L�ի��·��X�հ���"���Ű��r���F�������y��|����pu����[g���`cc��(
��v���H ��ʊaL>�c��������-���r��b�`aVDOO2�4l�+�f�Z�(D�4�/ ?❈�����LGſ�����8ݳ�p�D"9�uQ����n�8t�:�6���!���@�T�0���l6�H$'�y�^T�U�|�<�V>�n��%U(F�\���,ʌn�Z���r���ƆB!h��f�E��NUUT*�j5x�8��� ���H&S �����GDtE$I�z�
�x�t2����������'�x-F@4�������߿��nii��k)#���~����m�\��ϟ?��^�&G�lll��r�}]�u�1dʒ�b��a���>�#�-Q��,ݪYvޔJE�z�������u���0%""�G��DDD7$I�o4M۞uDD�A�Xv�}l���D>��0����*�N���Ӌ].��-��TUE$5��x<\�=C�Zʹ�JE��~
����U*�p�ܦ���� h4��N���`�|>�n���Y�o��$!
�P��n�X�NDsL@,���/_#�H��3���9??���>���r��([�����l���������6����y���(+�9�hKK+�1�^��� xl�׋���1�b�S�-���i�l��n�������?�p8<�4<]�qqqf�IE���i�?�0-""�G��DDD7$�bIӴ�:�<�� @�aX�k��Q��8�fʺ�.R)�)�v�J\Kl�N��H$jx��p8�����pg4MC��A<�0�s8E�'�=t��%<��d~ C�$��W�A��A.������x2�u�{*� �Н���ua�+�Ri�l�[�:��"vwߣR��3�~�����*$��yU���L�e�}�������b��3$"^�zm����� �nע�h}}��W�u�sʔ�Ad2ˆ1�?�p�)�%	Ít�����l#��_QU��DDDD7�w""��4�Tſ�����`ݳn��t:Q��H�h�`��FQF�x<����n7��[���!�0.������s<���~�Y����� :�6��J�>�.�y�{ �(���Y�NWt]G�^G�T��f���p�B�D"U��鰘����X,���H�o[�T����"��q�6�)�D�����{�=����ֶ�=�����}�~�oQV�s2�c��*NO?[��|>��Oo��,#��F�i[]}n�,VQ|�p�g~Dw �"2�%��'�R.�7`���R忰0%""�'��DDD� Iҿ�i��h""���nx0�v����Y�0e�^�T�0��p�T*Z���}x�^����dY�:�jaf�c�F�t�> ����%(
�A>d���\.ߠ�=�ݎj�bAv�X(����2*�K�\�[M
�e�H�x���������X[[/�N/�^G��j�pxx���/�2K��d2���L�l��v���=�����3�q�?��\��Yr8��~eXT��:��w�޳��Ʀ�����áE�'�݁����l�����( ��:�G!�=7<��$�j��,L����I`�;�-H��h���g�p59�Ncܡ� PU�F�����p8���3\Q�r�Q��0p��UZ�&R��ၗ��G�r������\C"�4<�E�@ �B �T6��e8���>���
M�O�(�h6p�=p87�7�ݓ�dYF�Ն�kSȖ��
b��|�
�T�օ�A''�p||�~�w�9�S�J���>Yq{��ûw����#������m:��^����Ȣ�h���-x�^Ø\.�b�`QF�����fS�TpqqnQF�+�YB02��qxx�!	Dw�H$'z�7��������f���~�(%""�'��DDD��iڮ  w���)��?`8���r#���0������J�c�N'-�(
$IB #</
����я)���h�H$j�p8 I'�?�~U����t:M�}>;���g��}��9t�]x�>�l���$!"�LA�$��mh݉�q�x�ka{�V�� 0����)�j5�9Kz*2�%<�b��n��w�gq�# �6�}�����h4���;�*�Bg)��ٳU�Eaoo�״���2�.u5���-�IElnnC�Ɨ�T*U�rY�"zzDQD&�l�G@�r�v�5�uA���5S"""z2X�NDDt;�,�QӴ�Y'BD ��ba!>�uY������-�j��Cx�fS�]h4����f6�Z�&��dY�t:1�n�=2+�v.��tB��@��A�۵(3�-]�Q.����L�  |݂�B�riAv�u��r9�F#x�>Â�q��S�4dYF��Bw"z�$IB:���/_!Oܺ�]U���a�z��m8��2�%���׮��9�����z	��o�c���3&�"^�zc�����'nk�P 0m:�����v��	��㟃��O�������.�� B���xr�,F����eY�#M��S"""z2X�NDDtK�(4M���΃��Z	�H�\nN��@���:�}�d���i��u�A��q_Z @��g���jUD�1Ӄ�p8�r��Uӏ�u�����5�������"w2���j"��AQF��nW�.�"� ��4z�.?S������XZZ���6��ح>瀫F苋s���Z�@�y�K�={����gŶ�m�{�{�Bz82�%�Ӌ�q_�|A>�g�����h4f�j�p||dQF ��ۦ�����c���m������z=|������d25�V�y7���oO�$��4�{�R"""zRX�NDDtK���N�?�Q#��DQ4��a���l689|�F�<<�����߅ź�.�~�a��$I�$	�j�����t]G�QG"�� �c�
S(�@�\�{<���?�y<^x�>\^�����t]G��D.��a��m
@A���G:�����h4��3͌�����3lnn#ݺ�]�T�r9���R�d'��������D��v;;�X��H��~lmmC�a��uZ���r�&�}]M���5�B���Wc���Y��p8l�}uv��fâ���&Q���,�^?P��?sA�TU�K xSFDDt,p'""���$IM���!"�N��T*Q_j��P*-�j>u:]��fS�]��n�V��d2e�`���V��x�F�F�"��a���,˨V�eFw�������k�v�qyɢ<2��W���E���7�O���F<�@4��i�v;��/��	x�b/^����ߺ�D�5
y���\.AU�{Δ�A����x<1Q|�uUܮ(,ndن7o�1ݐ5�����m6����m������,ʈ `ss�d�����}6�X�ŋ�\��������>G ��`0�P(4�4�B!gx� ��i���)=),p'""�Y�W4M�3�΃��*f�����cc\.7./�<p���h��mX��p8�j����,�l�)�Q��	��|l>��v����׸�������a�cQ�\��t��n��m�H���,�#SW���s�u^�������@4C<�� �v�,� �{'�"�������2����h��\.���=�JE~o�DDQ«W��7�^k4����EЏ���/_��������C�Ӷ$+/[��Ҳa�h4���.�M-����bS*��˱�`�</���c��T*��HtW�T
�Qc�����87�E��4���(%""�'��DDDw�p8�+��_�:"�k�^�����?QQ�\Z��|�t�H�҆���ͩ[k6�XXX0�`g�;0�j�,̌~�V�!��N�C(��P�<�J�dE�v��X�j��c���i�������z��$�V��,���X\���v���c4�s�D4o�v2�%lm�D<��n�����*����9��nF�e�~�v�ɜ�z��;�{D����J�L�NOO��� \7�Ȳ�u����ͦEY lnn��p�}]�u�q���֞>G��]���$IB&�t�R�Ѩ�^��蚦�� �.����X�NDDt���DQ��t]���-"�{�(
<<����n
�<�O��(��:�6�ݮ���7]�����'�� 
��'3��:�:�a�fQ
�Q,��b�XT*����������lC,��Z�ʢ����h�����z}�C�� �׋T*�H$
M���rs�L ���s��o A�n<��
��������kV��ݎ7o���o~ �j��;����Balll����5}�(+2���*"��aL����O�eD �D��,ƔJE��l�6�Á���ϵR��b�`aVDOS(6ـJ�
�<����%I:�u���0%""�'��DDDw$�򷚦��uDD���>���S�A�a�)MW��F:m<����r������^/��� �(�n����fi4a8"���l6��n��%�2��P�V`��&*��$	����:�C=��麎v��l6�~���c���@4C"��$I���,,%��$IB2����62�%x<�;MB������V+,8�s�\��o�~����=��="N�o޼5m����y�����`ss���A�u���p�mBV���2�޾��Ea#��-/� 0.������{�J�?�芦i��8���ccdY�{����"""zrX�NDDtG�$�h���:"�k���PN�sl���A.�5|�Fw�(
'|>���ݎn�Sܭ�l6�L� ��'�{�^4��㧰����m8����������lX�݇j�
M�
�Mc%I��B�V�~ς��i��n���e��t�t:�t`+�2��3�z�PU��D��?���g���B4�Sc �z]��~Ƈh4꼏�[�x<x���g?V,pxx���GDE�y�.��0�(w�7�<�ۯLg��'S[,�aq1cS(P,rz��I����-���Җz����3�"z�dY��b�NM���h�V��8���(
V�܉���HӴ�(�S�u��у�(#,,�Ǿ.��Z���Yͧv��T�l���S�-��*t]7-����(�,꘱Z��H$
��n
��j5����1i6P�p���(�������� �n��� �ϣZ�@�;MTn��x�dv��^���s�D��ɲ�x<���M,//���6SN��h���>~<F���5)�Z0ě7ߘ^O_;??���є������=Q����gK?�D����1�� ��������K����F^�O_*�F43�9>>� �{Gf�ƣP,���X�F���)=I,p'""��$�M�6f�ѵn�����I�n��l�¬擪*p8���ccl6;z�.��Y��j"5.��~��u�Ң���:�:��I���p8�r��C�G�1!����Xl� �Iw2qyy�R�t�Bw �$�@ ��i��躆^���HDO��P(���5��o"�M\@<��븼,�ÇC�������,����א�Ɏ���pr�i�Y�}[\� �1�6 �J���dDfl6^�2o}@�ݶ(+�Xl�q�A>�C�T�(��%67��qw�]|���¬���tz���3�@�u���6�ɲ�5M���EDD�$��������x�i�0�<��~*��}�f���i���Z��|j�[H���|>��'rY���"�H�T*��eE?g4���n� �VW�!�E���N��v��h46Q�q0��fC�V� ;z�e�J��|>UU�v{&.�y\.b��Ri8�N(�����r&��r��H�����tz��2�Ն�\.���}��y��̠���;�m�������gdF�)ass��s������w�4͢������0�j����'eD�UA�˗��5M���TU�0��tuO�2�����mn)%�+��n��CWZ�&�Պa��f��UU5""""S,p'""��������t]�ԓ��b�N�Tʰ@��p�P�Z�iSUv�~���KY�1��j5-̌�>\.�^��A����^y ��.DQD 4����p����,[�ݗ^��z��X,Q4l�����xQ�T��@w�i�:��,:�d���u�S�$�|~$�)$I8��}n� z�dYF<����/����`0Y�����z=�����p��%?�^��/ֱ�����B�5�X�=�c�p8���7��y��bg�{6�=�pϞ��躆����FeE�UcP<n�X��eQ.�,�h�mll��p�}}4�ÇC> ��h>�o�i<
�b�^o��(VE�[�DDD�d������H���j��|�y]�u��$��N��Z��h��H�ӆ��|>?r�t��Ԭ�l6�L&�iEA���Y�����}p�܆q����i��V+�F��$��A�ۍP(�J��(���v;(�V+n�ݧ3˲�@ �tz�P� ������E�h���X_�D4�����:*�
>~<§O�l6�Y@�FElmm�n����*��vQ�\N93�o�(�͛7��F pxx�z�nAVdF�d�y�ִI����e6m[I�$lo�2l�4��n�@ �Qk���3����Ft2�d�s��躎��3��7Y��M��w�"""z�X�NDDtOl6[IU�o�y�X��E:�hX�%�2�,����m�H�]�y�l1UU1���� ���j> �j�؂��p ��h4����eF�e4��H$j�{��P����*����CT*����p�=�2���t"�bq1�?�C�;�܈fO�B!��<���&���	�2    IDATn���\ @Q��9�#������f���oG&�W������Z_�@$5�;;��l��hϟ?G(2��v�8<��Tj�-/� 1����8�8�<�n�g��W��l$�.�k���y�n�LC%I�+��q5�=`�;�=QU��(�[���W;�MS�r����_-�v�Q,Y�k�V��d2e8	����X,p����6� \.��A��xP,����i��z��x<Q�A����%��!EQP.�
�`��M�m6P�70r3	�/M��j5��f�n7!�\.ם^��û�ư������Q�;���""��0��W����d2��kx�q�F������!*�
�h*\.޾�^�w��~��w�G�ݚrf4��"���M�j���-Ȉ&��������R���.��,f�ٱ����_Q챠�N�/^��o��9m!�'qx<�]CλR��^�;�uQ������DDD��������I��g5M[�uDD?��]Mq��@G�V�.�9u} 
���� I�P�T�J��j4H&S���N��~�N�����FC��}�bƓ�%IB @�Xd��#��*J�|>�a�5I���G��1<l"��^��r��|>EQ�t:'�4`��=�*v�nP��N4�("
cii�kQ{�^�ڇ�!r�,��q~~�N��k��?��o����(��n�ݻ߳���
C���6m����x���}Q����l�ͻ�\�\΢����ښ��E 8=��Z�fQF��ٳU��~Ø���F��Ft2�eá<�'..��$I��4M���DDD���
����ɲ�TU�ߚuDD?6���O��x���r�@d�v��D"Y������\.��b��@�4���  r����t �2�~�Ch���ۃr�dQft�t]C�T��n��7~#�5Q��� ���dH�JUU4d��V��<7��ű� ��� [@&��P(I�0��Ct�$!�`yy���E�{+j�j�����V�򚞦.[��W��1�V����(
�6#�Ӊ7o�1-B�4�߿C�׳(32����Xl�0f8`oo���,�r����i�42pxx�f5�l6lll^�U*��f�fE�ty�^��'���M7G����5M;�(%""�'��DDD�HU�CA���%�f4"O�}]Eh��F���Ӧ�:F#����ӂ �ᰳw������Q��p8qy�5�A�^���7����x ��s�X�R� ���A8�NT�U ,B����T*��r���O�5#�N'��3�D"�����M��p �H�ٳU��o ���v�j�C6{����rYt�𻇬���/^��N�V(pp����GJ�d�}������׎��^�C��x���e�^=<<@�͍qV������8�>��jY��|[^^A(2�9:����[H��C<����u�B�TD�;~c�(�UU�cS"""z�X|GDDt�dY�s��-�:"�����Fc��ǯA�z��岜Dd�N��h4j��p�=��kfF �j5�L��=:���m�N�ZE,�`:�2�����X�ݷz�����H$:Q!���C0B�R��q�5M��ih����s(�KPUN�s⩺�p8�BH�ӈ�_|^��)$ �Jcmm���G�r�&.����P(���G��|B�Q���(����B:=�#���3|�x4Ŭh�A�˗�o����s��sp��!�իWp:������|�bQNt���cm�aL����1??� I2���[�NOO,̊�����6�>e��g����$�3M��WS"""z�X�NDDt�$Ii���g��Oi�f85\%(��f�aaV�k0 �Ƹ\n
y�2�k���("0�Q(�9���4�F�D�`| �D�<�ȵ�m4�MD�щ��N'b�j��]��F���..��׫�un��^�m6�~?��82�%�!��v躆�pxo��Cg���D������M�RiA����Iᚮk�V�8;��Q�\�,g�;���7���뺎��#<?r/^�ca�� 4�[$����ɔa��������R3���e�|���!z=8�B&s������G. �'�@��=GW���FW�������ɢ�����܉��i;� �!�=KDL����B6�ml���)�V��z�_���<�Ӊv��C�h6��b���Oٗ$�,�Z�X��31y���D�H����8��=T*UD"щ&c˲�D�N�^ς����`�J����t�]� ��y�ӤA���B(F2�B"q�f\E�#6dѓ"���R��֞cm�9b�x��)L�Q�7p~~���C
yt:m�3�Lx�^�}�-�n�D�boo�riʙ�4�ӋX^^1���������9������+�念�#���H$���eØF��ϟ9-�
�(a{�%$i��Z���4}�{�L&M�|�J�T4��*�bOQ��������@��?�i��;���,���DI�0�j�,�j~u�]�)^^��|΢�蚮��t�H$ ��|>4u��}뒣�:��D��%�(�T*�8�����,#�6o]E��EA�մ C����K�r	_?��{/v�;|>?������u��p��wzTA���C<����3�x��D"�@  �}|C���h4���8Ǉ��]��j�}C3�-���7]� W�U;;ߣ�`��c
����ez���*vv������n��0�V����E�5A�����:��`��Z,�N/�-89��v�ϭ��$I�d���Y�S��:����%I�g���}�"""�,p'""�Y�۪���Y�AD�S�N�d�4~ڭ��E6��YO�p8����3���f�����n[�W!v�>�� J@0B�P�����!��k��+ ���p��(��W��æ(
J�"|>��F�k�  ��n��V�Z�!�x�����T*"�ˢ��BE8��)0�����|����,!
�PX?���C� ������X^^���:R�E�Ba�\�x� ?-j�f/�j59	�����x�>��~��»w�ss�#�v����[�i�Wt��ﱙ�I��H��g�h����(�bQVt-�H���jJ=�(��v�p�m��m0�Ç�3k��G	�+�v�ʥa��n�OE��""�{�w""�)PUuO�?�k�聹.\
��ccdYF��C�Âj+�Zm��)�B�߇\.�³h4���l�,�f��R�X��T*��p8�qn��(�^�Y�M��i(�J_��&��Ϗ`0�j���Ez4MC��F�TD6�E�������� ��t""O �YB4���$�PU����,�
��H$��rUțJ�
������ ��?����f/ptĢvzx$I���K����\.cw�=e4��h�dن�o�5���O�>�X,X�M��t����E�ﯓ�T�|�`5Q���k�g=��coo��I&S���1����l����,.f����)�
����(vG��haJDDDs�EwDDDS"��iZf�y������0�ۃ\.gaV�KQ���)�$C�TNc�]���v���|>Z�'$>���R�baa��� � ���$<�Z���pd��N�q4����E�4t:�&F�Z-h���1���v�~���3H$����_����sZ"���p�t��kX[{���8����EUUT*�8;������s,j���r�͛on4Y���GGG�.��	��ׯ_����
y|��a����/_��vF�ZM}�('����ΘaL>�C�X�(��&��^�f�����8<<���{�p8�JM�@9�t]���4m���$I���i��´����܉���D�喪�q�y����E�`hl��fC���az(MW��B*�6�����P(�i,��Z�׃����5��(���:���ټ��oV$
��h�Y����-4�D"Q�i����x<��h�v�eA�D7��:z�.*�K\\\�V�b4�n���Y���z�D�L�����H$
����]�9ђ&�t����,6�=���,���ZX�U��}ѽ�=m�� y8�p�	�8A� �'�d&���ü��@���<$�80@ g����$R$k�O�g�E]]�Ꜣ�x�H~?� ]�W�/�DV�9���H$�T*���9<}���3���p8nj`��C>�Û7�qtt�|>�f���m4�&&&�����=T���88x��󷷜�찴�l�| �j{{�6$�����A:�6�1;;���z6��k���k��5M�����$�L"�2��9=}�Z�jS"��/�H��7��MW����VQ�=]�Om�DDD����"""�(�]]׹ߍ�Ǝ,���/���dcEQ���1��677���G�5��%�{��,�����r=|.��˗{6��a��q���[���}|��o�j�lHE����`}}�rj�r�,��Hw���A4E4:�p8|k���h�Ei@Q4�ʻ��4�P	���P�������~��1>�0�j5T*e��%nj�;eff�?ư����>vww��wO��?��ܼe]���o�ͻ+4.�^/~��_X�}��5NO���~dqqɲ��Ϗ�~��߃���uUU�_�9�}A���ﶵ����7(���.������"""�,�{�����'E�/t]��Q� "�����d.133;����#�@�l>������H��L/,�R)d2�h48e�n����� �뛦u�d�R�B��dd�P(���e����������[Nѻ��6���X[[3�X�dr^���;�v;�����tڸ�����DQD(B4:�h4
�wp�ȗ$IB�0B������:���������0l�E���t���������B��gܖn��r��r��J�Mc�-�$cyy�Xl��4�
vv�����}�H$�jn�4;;/��>fA���es��4pv�!�����19�2���{܆a�X,n�� �ln'�������}��͈���?���w""�[�r��z����F����S'��_�˦7���:���[S=l���>]4��V�x��;��ǖ������7���M�cfee�DҲ��h���︊��O�.ZN��P����ގ�,�q�r��DG���t�o ����h�Zh�[h�Zh6���̛��Ix<x�>x�^x<^x�W��6A�EUUT�UT�T*�Z�QG"�l>�kk�x<C?�X,���=�o�'��677-
����m#C�l��u���7h6��5
[[�,@���¦D���?C �uM��_�9�}A��s�F'F�N��jx��ĴF�忢���������Uh""�{����� t�}7�G��2�KLMM�	��èV�����%��)��E�p�X�"'�����1"�\.���Á�O����mc2�rp�n����� ������m'�u�a��� ���ɓ'CMv:����
��Gll�;��� �� ��  �^/��Ȼ_a8�3����j����t��t�h�;�t�?�3�Yn�$I�x<p�=p��������� �όM�P��P�VP�V�(
_��^H$X\\�$IC>����)޼ynƸ�8��^������c���cnnβ���Wln�x<n���j���\ڔ��Ѩis;pu�����Q��	 P��M�.�b���DDD���DDD�L��?SU�_u"�Oy���t��&����mbNN����̴na�	��������x��%��̟�X,�D"�|>gS2���:vww���?��e~�0��ӧ�8<<�)ݶ��(�������0_O~�D"88x�u�t�ZW�үm��}���~�F��\x�P�Ƨ�k��v��n��n��^��N��^��n����(�p:]p�~���t��v�����ðTUE�^C�VC�VE�^gC;�+�(����C��4/_����=�v����l���<�9�DQ�����z����s�RчAģG�u''G|�a��Y�C!����۷6�!z��0Dq�C������5�(�)���.6��2I����D4���.r�&'Sk"�(��������J��R�����kB�n7��gpvvjc2�V�Vpyy�tzʴ���E�jUt�]����^�����x��k��T*�N���{�^��o~������U�bq�|>���BQ�[NHd��@Q��MVn��P�P�`�t���$I0������������������~�^��B��;�/�"$I������N���v���Q\��N��Z������f�N�����rcuu�r�ЇZ�vw��j�n1�I�e��ouЬT*���؆TtSss����O~8����ј�����1�)�J(��'�җ�
�.�f3��xM��K�D�s���k�u�k� �c��=X�_����E���{�9��>������%a�ǃb����mS=l�?���AO��4����x�gDDQ������J/^<�)+ccc��{��˗���6�"���G�cffv��躎W�N8q�Yv 
"" ����2����/M�`����~�U�a�д&�]�~����m� \5�_�$���	� Y����e	��x��I�!��P�[w��ih4h4�h4��j|_KF,����P���JE�|�ϭ2�� ����D$��m4�x���;{@�>�x��k�kj ptt���#�t:�{��KH�����a��o~�D6���B4�u�0��_�:������7�Á��u��,����	j��C�DQ��>�"""�l��NDDdQ����u�9��>��n�P( �H���b��|h6�6&{���6.//0==3�F�$<z��6&�k����`Ϟ}���H�T
�Lƾpd�Z����%VVV-k������P�p��}a^�:A��`qqy��QQ���SA����=U�T*�T*��;�����= �?�P(Y��M� ��xN��0�ۭw���5(��)���|�!;�0pvv�7oހ�塚���6�����s������F�J����z�h��� ..���n�@ `�� �|���D_X4:���!i��z�nZ#I�?�uݴ����~:ɺ����~*QOt]�wG���h�v��tzʴ��p�P�۔���:&'S?���1�߇r��i�#��v!�2���i]8A����1s}`'6o*�X�r	�^ώhd�f��r��h4:�U�ߏX,�Z��~�3�C�i����*��޾}�B!�Z��v�UU!��&�����P��Q*qyy���78>>�����"�:_O�Ar�\���D"��1������Y��o� �N[���}<�=�]6y��'O�"�0�QU���y@aD�~?a6���g�.ؤh���ex�^�
/_��37�633���C�Tʦ��@��?�4�hS$""���DDD6�u�\���0ר�}J��C 4�����P*ِb�С�:&&�n�
��|lx�Z��X,��9�FE�!d�Yp��x�ժp��&�E1
y6&�3�^�|~ �g��8LN�����(�[NH4���>Z�&��
��<..�qqq�r�EQ��v��:$I2=�Gw��ih6�����^��͛7�岨T�h6~v 011���-x<f�|?�(
�?������4��Y�麆���h6R�ME�x��e���e�ݞ��5����NNNP�UmJD�@ OLk
�"�}a~��F-���s�ϲ�(�UU�##=X��@DDdY��麾>�DD�t:m�R�ĜN���HQ�b1��i�ˍv��~5��0��u�R)��.�� �Z�ؘ��Q.����-���,�����u�|�("2��pMLL��v�Q�V`<�BtM�ut�4u�J%d��}{���s����{�.�eפ�1UU�h4P��Q(�qqq�ׯ_�իW�d.Q,Q������H�A����'O!��ߎ�f3������{(�Hbii	fӤ��ϙ��{�T��q9NlnnY�+��x���M��c�D�ӳ�5�V��6%" XZZ�<\~p��C�D_��dz��]����Źi�(���a��M����4�b�-    IDAT!""��(���m�9�����TʈD�kb�� N���a8>>���3ӺǏ��T*��hD����S��͛���΢R���}�\7�lm=C04��x<X_��������1�^]M�[^^�,;�z��d
�p��{��9����u����#A�����������ß�B�v��n��v��N��v��N�?��:�Dw������*�~�MA�u��G�d.o1���D��+�jn���c���E�eii�tp�再ӣ#�"=Z��;>>�ae�B!D���;@�T�ug�/L�$���QǸ3�9`�i�?�!
a��(DDD�ň���u=>�DD��!|��צ5�r	��/lJD ����X,fZ���k����'�A���?���7��v����@U9�q�8|��φ�fT�V�����ې���r�����`p�i��U����)NO߰A��s8p�\p���~�������d�D�u�z=t�]t��z=t:�z]t�?�����drO�.ZNw�P�����7s�S�`h��� pvvʩ�clzzO,���v�q����1?�ȴ�X,`wwǦD [[�GLk~��o�h�mJD�0LL�03c�т~pp��v�=��$�j�6o_"""����o���l$����:� �z�r	�����ht�P�Z��d���1��(DQX3;;�l6�n�cc2�f:��v��´i��raii�7Q�P�����s|���p8̧�����aww����P������G�}P���#
���}t�l%�R��>��>EX#�2�N'ǻ_���o�C�,ːedY�]���i*TU�������{�����z��՟��>�,cqq	�x�F���r8::���{���cccs���B!�ׯ_ې�>���ãG�-��,��G��rY~�3�^�ؔ�����V���b���D�`bb���N�c�� �$�S�o'""��ݻ�ODDt�% �F���L ��_�ܴ�R��ŋ�mJD �����|>���=�ѧ�Ri,..Y��D&��!�T(���3�%ײ�^ڐ�Feb"������3"TU���!�y��'g�$�kx��%I2$I�(�E�$AȲ��w ������q㢦i0�o��u�~u#\U��������]��5�����p8����\����W�緘�F���⫯��<@ �j��Ϲ%jL������9|>�i]��Ʒ�~M�������"�H�ּ}{�w�mm}�p8lZ��1=�JD7�v{���2�wF&s�\.;�� �a� 4�KEDD��q�;���$�i��]pD4��J�"&&bk"���0�UNq����$��p:�O$��d2�V+6&�e2��D"�S��V���jٔ��U�հ�����u��\���TU��ɱM��n�R�|����!�Y�����h4���CNc%S��A�4n\ ���z����n2S��naww�&��+�˅�ͭ���E���6��������v�0�����G(
[6���=���ڔ�  �Z6�
y6��No��J�l�uI�^����v"""Y��#""�/��p�4M��Q� "2�l6�N�av����"��j�\O���< �P(�L&�0lJF�T*H&���EQD(B6���jܴZ-t:�w�o�J�`�a�V���l�i*��dY�� �~?b�8��:z��-&$""�Q�z����z�L9|s{>����6��c�[[���x-k��6^���~߆d�9��	<y�Բ�͛����6$�O�p8�u��G���6�" X^^���6�0���ǟ�D_� ���jK%ͦ�B��u\���J��_������w"""�i��+A�7��EDd�~���o:���v�^����ؘ�aS�&&&��k�t]g��麎FCA29i:��tAET*��?��M��"��t�D��*�$���@�\F�QG$�$wI��p �JA�$T�5�@���J����nѰ�c������_���{L%lnn��X�v�]<�;�1�Ӊ��-����Z��6��O���E"a�MOQڔ���"��s�5�|���6%"z8���P�5�J.�E�=x۪ ��i W�وG�����ה$��CY9=}�F���G���w��[V���ݨт��Z����u333�D"6$��qqq>���'O�X�L���\.��o�r�4�cA���,~�������b:"""�mn�[[ϰ��4�7 h4����� �a�}&"����,k��>^�xΡcniiN�ӴFUU�|�σ+#�v�-�����<tl���yӯ����7�d!zh��>���U�I���UDDD6�w""��$I�u���:��~����op3���F�QG�ݶ1����v�v{L�$A���\�I��Z�"1���D"���uG�jN��@ТR@,C�����{N�4��9���p8b���CN���)��i�DDDwP29���Mx��=���{{{���s�	����uLLX7�i��/���TlHF�kff���e���>����Ҋ�a�l6���s� �b1LOϚ��r9d��=���3C_�z�����0Y����i;6E"""�w��NDD4��#��јk6��S�B�^��٬^�ar2e:1���BQӵ�t�j���J/P�$^��<$��r�����ϴN��	��uNb| �:J�"B���T�k�  �"��V�AU��FDD4�N'VVV1;;g���c�n��۸��'�o� `yy��F'�б��c9%�F��`uuղ10�����nG4ţG�MkTU���6t]�)��ʚ�ge�0���UUmLE�0$I�QǸ32�Kt����
���4�_�1�æ:""��0dY�u]�ޛID4B����1��r��Hm3]סi��d�P(�L&�5�#��}�z=�b1�:��M�P�s��*���x�'v
��D"�z��&����#��@�e�VS��r��J�a���X<����&���5�lo�@���������e$�����a`����P-I����ey���ncww��\FHElllB��u''�<Tb�x<���iӚl6�\.kS"��evv�t8�@�T�}{fZ#�������`S$"""� ������|���5�DDVE�Ԕ�w���n*٥�P�F�r��Ȳ�0P��&�()���g9�;��Z����ڔ�n�X, ��v��	��x<�Z�f:����0P.��l6�D���x=�=
�Z�B�8����h\8,/�b~�f�A�����''��u�ҸX\\��dj������[ND?���
��i�a��y�C�#677�X,nZ�h4ptthS"�"`uu��ۉF$Y�l���%��5�I�����FDD4lp'""UU_����0CD4b������N�s:�h�N��Y��`r2ez� 
�P(���ۘ�>V�V�H$!�����f�\.�f�1e��"��	�i~�("��Z���㡅���j!���������8�ǃ��TU��4n1!#�Hbcc��ͦ���u�x�=���-%�q���"�驡j_�:����-'��jjj33��u�_�B���!��x���jzM0����A6K$��?3�K�!�%����p����[�{'�(�4M��l�DDDD`�;�ɲ������sYQ��w���)�6��zp:��kA�������u�� ��4�>�e>��7�Ƙ��(������0_�.�W�ܫ�
z��M	i�4MC.�E��C8�(�C=NELL��DQ��x(���h�N��W177w���a����|@?^����P���opvvzˉ�
�C4L�Z������*�^�My����dx��N� `uu��z�����ۅ�i6&#z��g,_��J�ӱ|�E����l�DDDDa�;�9��4M����ADdE�T�\.�Fj�Ӊv��f�ic2��j��L�6`x<�Z-�Z|nF���@��a�:��]�-W���躆r��x<a:��a�{�\b���(��9���M�r��H��E�Z�q{!����T*���M���=��lb{�9�yNr~H?^j�7 \\��ի�[ND?�,���zfy�����ŋ�PUզd�)�x��s�5�~��;ܐg���I�RiӚ��n@ �%�D��[��|>gy?�0�? �ؓ����>�w""��4�"I��1�W�h�)���)�)�@ ��%�yv1�~�Xܴ.
#����ވU�5�BAx<Ӻp8�j��n�cS2�)UUQ*��!I�M�$!��T*���QU��4�H$An���A�X,�F��^�{�I���.�ǃ��LMM�y���~~�{{{|�~`��Y6�^�f3��}G���"Y�����hؐ��$	�뛖�͏��h�mJE�����u���ۉn� ����&�������~�$I'�a�c#�G�Ά��h�GRӴ�2�DDV4M���D08x��,�PU�:o ٩�T��vn��$	�(�R)ۘ�>�R� ��4�� "�(r�,%���&��I�V7����9���Q����� \.�Џs:�H�Rp�\�V�<<FDD�	����Y���[>�X�����6r�,�m�a���ţG����f�888��D�%LO�`zzƲ�����6$"3�/ ����j5��ٔ��MO� O�֜��E�X�)���,����:�Ţi�$I����fS$"""�6����i.�<��hL�0�}�d��)�lʵ��4�J�-&�Q*���lLF�4��@29i�|ɲ�@ �|>gc:�)U�R)����Q,��������f��4�P��{��$I�Z-t:�[�IDD��!lnn"�H��5�J&s���nZz���g���d��B!���}� ���X]]��YP�Uqp�ҦT4�����Ҋ��evv����ڗ�dف��u�m(��aoo�׌�n���4\.��c��l��:� ��� �?����F��DDD�דe�_�u�|���4�$!
��n�V+v�"\5O^=7�Wj� �ߏl6kc2��N�!&��ֹ�躎Z�fG,�L��U�{"�4��\\��b(��46�?4�z�r	�`N�s��ɲ�dr��z��܉��>�,;���S<}���� �n�������nUy�n�ܾ���'w�,���z��aZ������sR9���p�͛7���rP�<z����۷g(�K6%"zX'��gn|x��4oߞ��_�e�׺��c�'�����hH��w
��h�]O
7�T��eـg�Z��d2	Y�ָ\n��=4�ѧ�j5�Ax<ӺH$�z���)��S�׻Q�{<G�Tb�������f>c�;����J���:�?ǉ����LNbcc��a��_{������v�ns��C433;ts{�X`s�����`0hQe`ww��ؒ����F*�6��v���������n7���'���}����08��6$	�QǸ3*�
j��i�,�_�4�o!""16��]׿���f"�t]�a�F�kA�$�(��6&#�0��u��/	��<�0&���% "�(����1���P�Uo0�=�R��&��^��P������6?��!Q�N`b"�f��n�{�)����6�Ϗ��uLOO����fS������%���Y<~�0Tm�\fc�2;;���)˺��Sd���ˍ��u��ه�/ya�<yj�X���	�un'$�� `nn���u���s����_E����ic$"""��p���ƃ!����>�"�k4�w���q���(���6&�V��n*�w`�(��z�\�<t]G��@29i:�J�$��>gw@��E�VC<�z�{�\���JUU�rYt:��a����N'R�<j�t�������I����y����� p��������v�E�z��1��U[.������cwD(��6\Mw=<<�)�YYY���7��T�x���M�������"̶�t:m � ��
�11u�;������´F���E���ɦHDDDd��DDDcB��=]���Q� "�U�#��.��|��\ �F�T��f���E��F�ٴ1}J�ہ��DoE  ��AP�VlJF������.I2���2���fSA.�������c�~?R���3DDD��D[���Y6�~�V�bg�
�؈�p=z���sC��jU6��!N�[[[[Ԯ�smo?��1�H$-�u]���nG����! pxx�f����n���4\.רc��B�rۇ���[���l�DDDD&��NDD4&t]ψ����0�HD4&��b�	8��/�z�^�jUt:�zg��z�HĴ.#���F���k���z���Ba�Z-�Z<�0����x<a�X%I��*�2z���q�~�4�B�V�P�F��EQD4:�h4Ei��=H^�++k����l^����8::���>pO�<����P��Z��/�}G����M�I���������^�~�R�}�v��x��iM�Q��ɱM���˅��QǸS��NM߻���VU����HDDDd��DDDcD��i]�9�DD��v;H&'Mk�^�ٌM��Z�^�Ą�I��t:Q,mLF�T*e$I�f�ht�R��7w@�݆�(���C5�'	T�6'?p�V�lN�~�U�͏�\n�Ri�\.���:�������e�/`ii��Ə/���y�Z�v�������tzj��j�j�?��O�',�^�~�\.kC"�����`0dZ�l*88xiS"������胃}>!�E�����Z�^G�X0��$�Ot]��m�DDDD��NDD4Ft]��A�# 7۟LD4"�v�Pش���r��l��j٘���)I�Tڴ�����Ѩ��nۘ�>E�u��uLNN�>g�("�"��r���n�Q���' ��i�(^Mr��j�v�6%�q��:J�"��*� �N�Џ�@ ��DQD�^�a�����hT$�����@8�<P��v���/�-�8��'����J���gs�ݓLNZN��J����C��p8���'�5�a`gg���G �H`jjڴ�\.���ԦDD�(�������H?�d.M�����/��<""�1�w""��ғe�_�u=9� DD�j6��i���	�����/ z�$IB(d>�*
#�Ͱr�z]h��h4jZ�p8����ϛO�����tP���."�H�^�s���� ��D��G(��MKQ��H$����j5o1)������בNOA�nv��0t������.bӻ��eLN���/����y���wH ��چ�!�n��/����1 �677!�Ӻ�󷜶?� `mm���c`oo��nQ$E$b~�~��*޾=3��e�W����"���NDD4fdY�k���F���hX�^^�>�o`���@�ۅ�4lLF P�ՐH$Mo:ɲQQ��mLF���u�|��S ��z!W�i�u�7kr���lr���:��,�N�����v8����P�>�����x<X\\���7�pr�Z�`gg�|�|	� `ee��p�FJ�"��v��~�8lm=�hĽ:�����v��^�����F'Lk:���w��|����L�����rvBt�ff�,_���R�zݴ��p�]Mӎl�DDDDC`�;ј�4m[�?2Cu"�a)J����4�`0���K�x��ah6�it�`�J�k��D�\��D̲i'��jr����vP�Vn0�=EQ�n�mJH�L�4�E�j5����t�=H���x<����uN�$"��C�$���cee�Ƈ���MIGGG899F�߿��t׈�����b������L{��������ڣ�C�JER��@ ���%ˉ�{{;�2�$auu�t{�����݁��6&#zX|>���g����Tu��%Q���;6F"""�!�����hI��]חG���hX����t"��$	���V�i�u:��n����� 2� ް5�0P.��LN��4�ht�b��:wD��E�RA<�|nAD"�@��A��ؔ��]��A6��aC��?&���#�J�:��&-""g� bjj
kk�F'n��w�����-��v�hp�]�e��D�C�
y����}����d����\o޼�!Y�:��	��eZ��fp~~nS*����#�����oQ,lJD�0�RS�x<��qg�Z��
�    IDAT-�rY�Y��G]��W�"ѐ��NDD4��w����Q� "��F��t:m:�8"��@�85�n�Z��$dy����	�0xaL��
EQ�H$MyDQD$A>����6&�����P���'�hr�ši��]z8�V
y��x��=���F��)�j�Ҽ��DDD�/�H`mm�d��=ӧT*��l#�ϱ1��s:���|fz@�C�|/_�����H$���Ĳ�^�coo�����<���������#�t:���jz�WUU�����!�E�,cff��?�l6�v�|����UUy񕈈h̰����hi�V�$���a�?��hL�AGֈ�QQ.�mLF�����v�'L�B�
N�N L�� ��p����P�����^��R��n����'ע�($IB�R�!���"�ϡ^�����t���,#�#�H����b�;�^(�����g�p8n��v����C�~}��5�#n�[[�������d288x	n9�[|>?666 ��p���d/^|UUmJFf�^/VVV-6��(�p6
O�Lk޼y�j��-�nS<���]�y����0�$I�z��?�1��DDDc��pD4M��Q� "��F���ɔ��@ �b��F�h�Z����z���@ ٬��N�O�V���l��z��:�lJF?U��G�\B,7��y-
��p�\��b��N��L��n�`��Sn����(�����-%%""������E,,<�����5M�۷g���C���G�1�׋����v{���d.qxx6��-�����3˃��a`ww�&x�kk�x̿?K�޼ymS&�����ӧK���.7^�`nn���=T�J����,�����aS$"""���!""S���� �|��1��ab"6�Fx<^�rl��Z��T*e�N��rAU�h4��s\\5A��p�ߤ�D�h4h��6%�����T*����Q*�lHGw��4��\B����v�ܘ�L!�Ѩs�%���raa�	����?��@.����6J���w������������-��/O����PSmON��m�LMM#�N�֨�����4ͦT����x<^Ӛ��#(JæDDS(B,u�;���-z�������4������܉��Ɨ*��_�u}f�A��n��T��Mq=�pGD�4��jz ��0
�T���ǁa�V+���4=� ���@�X�sw����b�����e�����G�Td�]�Q�TP(��x,� ~���E:=�ӉfSa	�
�Ӊ��GX^^E0���,�j����.//�zE��D���5�aR x��5^�~u˩�6<~���ɔe].��s<F<VW�-�u\5O�jU�Rчb�8fg�Lk��&��mJD�pMO���r�:Ɲ��uqqqaZ#����������n��DDDcL�]���Q� "��^��D"iZ��\ڔ�>�(�BaӦGA9i���}4�-$	 ��DQD$E>�������DUU
yD"ѡ&Kz�^�Ba�E�g�]�~�|�z~`艥�A@ ���\.76�ї�p80;;���U�Ñ�jl�v�8>>��ɱ�DFz�&&bX[ۀ$w;���oߞ�r*���$�X�)������7,��jUnUQ���Y6?�p��v˦TD�����g��D>�G����H�􇺮�&јb�;��u�T���0���]$"�V��P(dz���p@UU��u�ѵz��T*m�L�r��i������L�݂ �æu��P�\ܮzwh��B!�P(��mY�v��DQ,x���t:�d.����n�v����T�,CQ�{#"��"����cee�H�rZ裡jo޼�˗{P��-���"������P������K\^��]
����nyXFU�x��9�}���s�S�u]������R7
33����5�r	��o�	D�MN����F��0gg��װDQ��4�?�1�܉��Ɯ,�S���r�9��n��P�N�7P�Ad�6ʍ���0�HԴ.
�T*�F��Vk�z��un�.��RѦd�%躎|>�@����9��LL�P*��i�	�j4긼�����7n*�P���N'�Ή�DDdM�$LO�`mm���CG6����*�
�/����9<}�8�v ]װ���B�`C2���n7���A�e�:�0����F�cƅ����ʪ���7�Q,��(8�N�����n_o�!��E	ss��>����k(�J�5�$�����ܦHDDD���NDD4�t]�A�O�|_3���}8�N��5�(B�$����v��uD"�Iт  !�͂���G�\B<���a�"��@UU4ܔp���B!����oY�p8�H$Q�V��q!f��2�  ���!Q�NOA�e4T#"�O���}��l�1P(����\.��2%�>]����P���b{����-'�� I�����m�����W��6��a����M��e�z��/mJE{��)���i���9r��M���X,�P�|�'����9z��������� pz�c�;���ɲ�7t]7��ID4���:��Dq�G�?�b���#R�U19�2m6q:� �j�jW,���:��
�ɤe�P$E�QG�ݶ)})�R�,[�P��;��$E�sM�t]G�RA�P�����ע��DwQ�l*l:$"" �,˘�����b��mlJ���v�o !2#IVWאLNU���������}G	����u�B֟���<NN�mHEÚ��D"iZ��:��_�z���~,..�l�����ρD6�����VB?��z��xkZ#������kS$"""�Llp'""�ǹ�i�ƨsݔ��0�ht`� �z���5"��B�4D��u�P�r�t�	٫��CQ$I�	̂  ��T*qe�T����:"��?G����D"�^�Ea�Y���(�(���x��?EE��LMM��t��lB�8����!r8������&&& I�w�Ѩ���}�����+��p`ccs��� ��t����h�����n���3(J;;;0n�~��˫���NN���q�VW�,�#����V�0��
���G�N��sh6�Q�����]�DDD4rlp'""�4M;E���u"��j4��p8k�n�M�V��dt��h �66
��P(�l6��c��n�;�`��!�"��	��9Nֺ�����>&&�0��\}�NL� I*��=�������P^���掛E�`��\.Z�&��=.��=���
"��gOlo��8::���1:��NI�������W���CշZ-<����a��)<~�`Y��u����PU��(bcc���F�V��ѡM��c�D�ӳ�5�V��6%"z�fff�t������٩�5pQ����6�"""���w""�;B��'��5�DD����X���d.�<="�Z�Tڴ��p@E6͎�z��˅@ `Z'�2�� ��<���F��v��X,f9�����v{8�n��n!���I��  bjj��V��w���)�ۍ��GX^^A(� |^c{����W'8<<@�ɉ�4�`0�����r���h4������z���nK(��ښ�g"]����R3�=��B�i����`�����ȲlZ����v�mS*����� ��u�;�V�Z^u8���ijS$"""�	��NDDtG��� �CX��$"C�v�`�w`�,;�i�����蚪��&D�L�B� ��*�]N�'�r�}C����ˍR�hS2����&Ey��n�@���Q*y��n��=�v���g��eA���155�χv��f2"�{����ɓ�X\\B0��ݧ��m����� �F����.�c}}Ӳ	�Z�\���n����n���A������=T*eRѰ���,_3���8Xa�fg�,!�E���ڔ��aK������B�������� ��i� ��"""���NDDtw�dY�C]�ͯ.�)Ei ��2�����f�i���蚢4," ��0��f�L�TB<�lD������mJF_R��B�RA,�$Y_��x<����T*�g+�X�����%Z�&�~�g5�|>��)D"Q��}�ۜ�IDt�B!<}��'O����vc{��g��b���4�?g�}_2"wo�;W���F �P��Z�	D��a����h��\p7h��F�0�@�������t��=c�#N�����U�W>'��8����T�]o؏*gy����۷����E���v����1���v�k���vv�aF��Q�H����x<����7��8w uJ%,--۞O
y:��~��vcnn�rwG�4�����BD�$�_|���Z-���Z�Ȳ��aǡHDDD����NDD4@dY������AD�%��6EA(�l�(�P�ӥ{�X,bx8Q���,+�$	�<����0P(�J�-oF@,E�Ze��R�2�,b�XG�.�����'h���k8;�����F��]$��RH�R �jU.�""�s�  ����,&'}��V���o�����r��� �"�=Ɠ'O��&��޽e��ϟ/Y^O�����wz�l
�X̲F�4ll�qavMO� Z֜�� ��v(��644��g����j��e��(C��#�"�Wb�;� �u}S���4MW��}�r����˩Á@ �|�M�=��:TU�ݎ8
�R)��h8��:�n�Q�V14����# O�6�4MC&s�p8��m[/�2��R�T�h6�$���^��讪*�~?dY��?GQ�bq�@E��uNT%"�3�,cttss��x�s>Nl���ac;}1Q�07����ю�M���ޮ�O�SS���+�J����{L��D���������E�Tr ��P(�gϦ,k�m��[<w#r� ��|���t�4M����=JŜ�i�`,"""�J<"""0�,?3�E�s}	�0��:��E� �ߏ���r���jUA���p���0M���'�f��!�z��옐H$��f���2��W��|������("�J��n�R�8���'�Jggg��k���P�/[+I��(FG����P���n��8/݆�����$fg��'�x1ps\���[Nl���r�����h�z�G��ckk�l��ɨ�&&&111i[�l6����s�>#�2���m?K�����JE�fnn�ǲ��� �r١DD[4���K?W,Q(X�8�(���u�w(�6��0�\�����KD�g��*�$\��7ù���u����IR���Ri�)1�,��v#��:��:Q���r�Zoc+I2b����8�k@���l6EQl�o�fT<���F>o}Ӈ��ǉ��z^�.חM��@ ����h���i���a�HO�<���4��DQ��?�V���� �(��ll�������~A' �����UN����!LOO��2���X__C�������,��eM�����:t]w(�R*���ؘeM�Z����C��h||���	����S˝JA0t]�� 8Y���h������h�4dY��0�{���K��u��i˚P(���s6C�ah6JY�4�j\��o
�<B�0�^�e����q}}��� ��s&����:�`0�`0�|>������:..�Q,�v{l�w>O���C:�F*��(J��k�7JD�%�(bh(���9��O���C�|�B�Z���x~@w"�Lbqq���b��VWW�hԻ���-�`a�9�n�����-�JEGrQ�R�&'�����p���$ϟ?�$YO�����"d"���~�Ӽ|�V��g�5�,��a��C����莰����h )�r����:їj6����|���e� �P(8��~�^������X�E�Qd2��
�e�Y��	ۉ?�>�����J��z��x<�Qs���E<���O��Z���.Q,�(.��y;�� �att��f�6�l��׋��I���ch(���!K�ptt�]��Ό��aff����b��kh�??�������Ҋ�r���ҁTt���K���\]]���w��_���SD�1˚L�'''%"���qx<�^�(WW���!�(��a|3#""0lp'""@�����7M��"X�J��#�M��P�\�rkI�b��T*Y��$'Q�xS����B!����ms���$�\T2���:��"�DG!.��T�J����δZ-\__!��A�$�|_>��3&���Q��躎F�qǉ���xSSSx�l
�p��巈L�D6����.޿ˉ�tgDQ���,&&&���D ��d���	]׻����rce�EGo...p|�ƁTt� `qq	^��bWUmass��5��������﵆a`kk����r�066�U�*=4�a�����;�J�t����8�����܉���,�#�a���9�����i�e�p��5� �����ӽb��:R��e�ǩ2�"��7���X,"�J�N?���4�J١t��V�|�X�rq�G�$ah(�V��Z��@Bz(TUE6���9���m�8Z�z�B:=Q�h4��FDd��raddss������?O�u���awwP��%%�������x<��c޿���=˦&�$ayy��]���vv��y�7�=F*������B��]?zG��狶S�ON�#��8�����G���{c���9�{�$��a�ȡHDDDt���NDD4���A�St:ʈ����e�����f�M�=�h4�(
B��e]$F�T��>��-�j5$�C��b�j��uN�d�v��W�Bmk,�$EA>�)�t�t]C�����TU����h���Ȳ�h4���q������DD?# ��ɓ����E,���]�f����	�����e9ɕ���������������.NOO���� 7ͶVC>��j��X�ap�c�	�ö������g��_3<<���Q˚V����m. "r�$I��|���tr�����A7���� b�;��j˲���1�� DD_�4M�Z-$�C�u�pܶ����"���6���./�\��F��v��x<nS) �H�X,���D�Af�����xt�(
����x��i��T�8;;C�Z����m� ��x�^$�C���B��d�%=Xn��Ӵ���1����n��V�x��{{�(<Χ���X\\�9��UU����|>��d䔙�9$�IۺV�����h�?��F�!�2��V�(�e]�V����7{HQ,,,B��[Evww8e��ACC)�3�s�ZWWֻ�ʲ���w�DDDDw��DDDL�m�0��^� "��z�P^�締�$	�,��u���r��tzزIF�ex�^d2ܾ�U*Ȳ�P�z*��4��٬���i"���4MD�ю����Ǒ��(L]�h�qyy�b�YV��z��	S�$��a���!��446�ѽ'�"�$�={���)D�_?�0���pp����#�E]59����E���Z����U6]�#�=��ؘm��iX__E��p ����,��e�a��X��r1}/MMM������C��HLN>�]xB?wqqf���$I��a�]�DDDԷxtDDD4��8E��5M���,DD_�R)cxxĲ�-�P�s�t��m躎X�z���G��d#L�*��z}��%IB<G&s]����T*�V�!�w�<�r�0<�F�^G�^w !=T�V��5��.a�&|>�W���8�}ddn��چ��w����?��O`vv�t^���Mk״6��ΰ�����s�f��!I��022�N����yln��s�I�����3�:�4����r��@*��T*���G�u��^�c�pϞM[�|\���DΉ���b��1P��6NN�[ֈ�x����v(u܉���$I�0��^� "���AED"V��A\^^8��~_�RF0������ �Ɛ�d8��O�r9�B��P�'�
"����9������r���MvECC)H��B��@Bz�4MC�P���)j�\.7<�W���$!
addCC)�\.4�-6j��r��H��1==�G�#
�ɔ�j���o�c{�    IDAT�����|>��I�:�ׇ���i�?uvv������d�X,�����v����A6�u ݖ������B�|>���C�Rѯ�p�\�uo�#����I��(J�c�L��jŲF����0��ϡHDDD�lp'""p�a�� �	��ND�\.#�JA�?!�f
��J���%uW�P@*��l�E�P����\.�D"a{���v���#��8�����Vq}}�H$����c��0�� ��<���L�D�^���ŧ�~����'+�r�`gll�h� ��h�4�o����(�H$�x��)������ru�n�4d��͛#T�.h$G��	,..���l!�i�8<<��wo���������Ro����܁Tt[� `qq^���v[���:w�뱱�q��i˚F����9(
ah(���4M����:� -]��y |C#""`l�#""|�,˿5�z_I"�>g�&�:R)�-�p���0���0P��l���ͳ�"'?�#�0��e�L�N���|�z���wO躎��+x<^������L&Q(�nsgr�����r��8��i�z��>`M���A<����8�� L�@�ټ��DDwA�b1<z����J���}�b h�Z8==���.//��G�����D��ۓ�����2��.'#'y�^,-�t4������oHE_���'5enoo�Z�:��>��ra~�����m��u�R ��Mt<��n�J�OC>GQ���0���P$"""�6��.��k��'��AD���� |��O~E���V�=�l6 �2B��e]$F�Tb�L��u�BCC)ۛ�~ .�b{��i��f30�h�}Ü�(H�Ө���M�2�R	��g(�ː$^��7z
� �ߏ��FFF��xa:���%'"��p������(�� �~��Ӽٽ�͛#�X,r�.9J�d��/`tt�w7���W���=�v������F�\.���Rї�#����=&?==����C��sfff-k���qr�ޡDD ������1pNOO���U�i�_��UDDD��DDD���iEY��U�0��BD������G,�m� J�"��{�T*"O��rYT	�F���~�P�v��J��Tj���t0p����P.�P����m9 7������bɁ�D?�h4��\����f���s�3�$!!����(�~?L�fAQ��ß�Z���!A����M�����9vvvpqq�F���y~ +++���*��bcc���'��`y��^�mm�R����#�)Y����l;��V�agg�i:��~M4œ'O-kt]����9ldd���E��f�i�pJ��U�0�+�"Q�����螐e9����:���x#�f����!\\�;�>�4M�J%[6F˲���m��X��D��"��_+�D��:����	�z�l�h̶AᆀH$�P(�|>Ǧ�	�0P�Vp~~�ig	����B;�$!|��>
��M��jYN#"������>���q�B!H�|'�a�f38::���
�t]��?�趆��������������1�I�����@ `[�h4���M�{W����G8l�h�0t����Mإ.ϟ/ٞ��A��w(���011�ջ�=4���;K*��7t]?t(u܉���	]�7EQ�LӴ�ߕ��ϕ�$�C�7_\.4Mc�m���mh��x<nY����i*>_��Z�ٱ5�^\ �X�F�Z�۱�!�v��W�z}=���!�L�X,��nw9!�穪�\.���3�Z-��.�\wsZt3�=�tz���p��0�ʉ�D�9AG066���YLLL"C�囹�9�{��vwwpuu�ݮ��Aĳg���ɳ��i����Mۉ�4xDQ���RGS��mkk�����FG�0>>n[wxx�|�ӽ699�drȲ�V�aooסDD����0�~��_�;�����w�;�����4��EDDD]�w""�{D�Q�4��DD_�D�VC:=lY�quu��s{�R� ��n��Fc(
�Q��J�"dY��@@"�@�ZA��p$u�a����avѰ� �(
��a��,�s�a�R�����L�ֆ�㹳ҏ���0FFF���!"Z����U"z�DQD,���8��g0::�P�n��UU���޼9���T*eN���s��X\\�m���z����U.`��A���b1�E� �����P�s!u�
C�����6���pt�����v{077o��hgg��&I2&'qz�-e�9�JE�I���0��L""""�6-�/>Aʦir�ss�JY�d2loo:��>GQ�|�ۭ�[�&^���Ӟ���̬�ঙt}}����x<����[5�]]]��`������CH��JA���T�0�J%�rYd2�PU���"�� �#�#�w�='�����
�|�l���C�A�?��/�rY���@׵.&�^���!�2���;x<�:UU����<&�ϟ/��xyy���D=�Nw��H?����V��rA�L�����=��7""���-��?e�d��݅r�����IC~��Z�z��d�K�a�V�!�J�j-�,�������r.�Z>��h*� H&����y}�4d�YD�Q(���� �$J�"�P_i�Z��r8;;E�^�(J�x<w6)Mx�^�bq���#�AQhZ������!�Ɠ'O�����$�~����1Q(���[������
�����G�czz��٭G�4q|���0M�<p=}�##��u�ibgg�BށT�����;������&j5N��dr��ַ�4������B�0Q19�����r��l6cY#���j��s(9��DDD��$I��a�;��ADtt]�a�[YG"Q\^^��L�5����p8bY�����:���s�l�H�v:�(�H&���l�g4����Kx�>�����(
��a��*��j�ݎi���j������9TU����}�6A���A4�����a�|>���V��I�D��$I������4&'!������*NOO������3�jU��P�q��x�|	�T�n�n���������y��1&&:������E�}n||��c�u�߿��Ņ�Ȋ,+X\\��I����RɡTD�Q"�D$b}��~����EQ����\1GDDt����V"""��(�7c��9��� �曗�u��g88�w(}� X^^�mr7Mkk�y#��I����A��V��ׯ��&�����<y��\J������>C�^0�;��x�'�L!��J��L�D�ZE>�C.�E�R���EDw���"�#O wu�b�^C&����w����F1;;��b�j[[h6y�p_���bjj��ڣ�C���t9}�P(����ϾR����U.����s}^�RƏ?�����A���.���&vw�-kdY��4m֡HDDD�Np'""��dYV��g{�����jUê�2�X,�����y�Ri�IQ�  ���꒓���i��H$�PŲV�e�b1d2�|N�r��j��X,�qS_ @"G�P��q�?�/M�P��qyy�L��v�r��݁��>�ۍH$�������CE��*�;����(���4�=�������v ��j��{��b�;�P_�?��������������}�c�T
333�da�۷�89y��P��dY��Ҋ���v[���4Ms(}N4�ӧ�,kL����&T��P*"�(���VK��������_Y��=]׷�DDDD�w""�{JŚa�^� "�+SS���i4����� �"�(���m���66�JE_���`e���n��J����U�ؾ��n��
�:~���������U��=�&��l6P(>}qa�s$IB(B4C$E0@�o��nR�5��ZW�.���(.���#�v��0�����N���z-�Hb~~���@gg�8<<p }���E$	�*���(�d��E	/_~��kYwzz���C�R�O�����~���麎���{>�(��������'��S�(N���m�sݕR��T*Y�?[�(
A@�Xp0��f�	A�D,�^�@�\r(}	MӐ�e144d;���vs��=����� �r�M�("�L��r�X,p�z?�잁�� �RG�}��,+�H&�0>>�x<��A��*_;DwH�$D�Q����'x�l
��0�����x7��M�����������i �bq,//��t��z����5�r�.&�^��b����nO��W���w }���I��Z� �w�����Dd�ɓ��ǭ'C7�Mloo�܂���0�ɡ^�8��5*��e��(������C�����A��NDDtA(��iW��h@�bq,..Y֘����jաT�y�����,�L����*J��C��K�!,/��6�@�\���t]w �B"���̜�£_�������{44�ˍx<�D"�H$�Q#��2M�r�R�r	�R�;e݂�(�������BM�Z�a�X, ��"��BUծ��D� �"=z���q���b6����.?��h4���;:&��r���`sm��#X^^���,�X__�����^����9[__�}��������u��b�&����n�<J�4� ��sɈ���)lp'""��dY�����^� "�Kss��tR�V��?�[p�\�����r�,�Z�^���,@$���RG��R	lr��<��v6��i�{��''' �>M�Mo�@��q��	�ϻ��l6P*�4���%�j5��n�~�r����=���!���P�#��!�˲���������Χ���7o�pvv��d���0���Q�����E���ի�x���o�yi�>}yy���]�R�O��LMM�:��)x��زF���IӴ��HDDD�06��c.�kNU��^� "�K����~EQ,뎎qzz�P*��D��d?��P(`cc�@<�����&�
ln��0�Q/���'O�btt�V�+
��݁�r���  � �#�9>�MU�O���r	�j��� ���@ �P(������& P��P(���P,y<K�F*����4DѾy��f����-���.&�~
����Ys{�V���k.��{����&�IE�&&&���˚v����� ꑧO��j8�88س[�oz���F��ADDD�܉���9I�t]��DDw)�Jcvvβ�0t����h4�"+������cۺ��7x�����k��i��̢�K�|[[�l����$fff!�rǏi�����E.��b2��p�\�Fc��o�ڸ�i�Ѩ�R��R��Z����bd� ���!"~����2wI�u��e�rY�rY4�MG�~�nS33����z\6�������P(���������:VW_����~�k7��������l�������\;���~���}��J��h�mw��eyUӴE"""�`�;�=�r��%UU�~�sݵ��e�b������VJD�:�f�7S��EN��p�7h���0x�>��/�n��K�8<<�a�]JF�[7��ÈFc���~���0>5��|��h48m��� �z}��B�7�T�V���P(�Q*����{+�bvv.���ǘ����789y��d�/� ��_t�x��h`m�5Z-�����(�mwj�����X���~����H$jY��尹��P""��Ǐ� ��:��y��-���e����k�V�s(� ܉�� Q�a��	�+�/_��vZ���..//JEVŅo�}	�ۺQ��n���$�1::�gϦ:��f3���bC�='�"����N��q�Z;;[v[���G�QD"Q���n2�Z�Z�j�Z�j���Y&zxE��@ �����W�� �j5Q(Q,P(䡪�<L��(�x��	���o��f����-T*�.%�~�����EQlk[�&VW_��~ ��|��K��UUU�z�=?����(���-kt]����%�����݉�~_�������5dQ��H;����z��DDD����/UU�۽�ADt�������3�M������������Wl'�U�U�~��ӾD'�ŏ2�vv���$�ILO�v4��#�0���1NNN�����x�^D"�_�\�^GB���I�{�Z�F����UDQ������Y3{/y|��*���ś��F���HD���|����.<��5����iZ��Q?��|X^~��qJ��������~'�"VV�A0��3Mkk�(��%#+.��}�[��탃}���9���~ir�1�Q�]��]\����ҲF�忥iڟ9����z��DDD�"B�4M��:DDE��/
�-�2�kloo9���LLL���'�uWW����q ݅�4��<��`����x0;;�p��}������v9�,�ǋh4�i�{'SR���*j���j����&��gdY�������������]��]�Q.�Q(�Q,P�Tz������ɓ'E���~J�5��������٨�x�>��t�ܮ�*��^�^�;������lG�o�ys����$�N,,,"�HX֔�%�~���B�n����}s�3(������JAZ�i� p>�=�#)""�B���QӴ?�u"�������/!�e����٬C����狈ǭo��45h=z���G�^^^`oo��z�	����q<~��V7�4MÛ7G��8�b:�A ���###
����:��Ѵ6��:��:��͛��F��v��U�#�����������tvd�e|�l6Q*�P.�P*Q����z�<fff��n�h�R���6w9x@�^��v��6�m�����k$��5::�gϦl���66�HD�H&�0?�`Yc^����E����D,�u����dpvvbY�(��m����3��������NDD�@x���F����'�{���ZUU���������(��ۗp���L���vɡd��?~���Ɏj���pp���D�/�������zo��L&���=���.%#<n������@_O��u�S�{�����f��V���>%�
�n<�/�o~��Χ=;�4MT����7_���u,���J�155}�ױi�8==����&�<�Ms���Is{kk�Q���v��,/��C6�M���<��,��~c�����޿�P*"�%Eqa~~������i����F���s7A�4� ��%#""�^���"��+MӾ�u"��&�"���;�|>˺��s���9����x�DѺ�BUU�������<y����r���"I�>}���[=��V����l6ӥdD�M�$�B!�Ba�!�A�\�^��a�h6[P�Z��}��v�͆�;"E��������������I�DU[(�+�T�(�˨T��u�ױ��������LG�i�T�����J�b��Q?�z}X^^騹]�4����R�8������·߾�m�6��?�y�#��sH�Җ5�Z�^��cg�G"��u��S,����Y����išHDDD�clp'""z@E�M����^� "�P(�/���i���:���3��V*����m]�\���k��@*�ϞMatt�����k��n����L&1==Y�o��L�����4N$��v�?5��|�n���7�v�v�U���7�V?�Z�t��`&�˲��/��EqAQ(������~o�iZ�J��W�J�!�:�Lajj����L����=�n�|7��v�����5T*e�����/�mk��vpyy�@*�D<����6U&^�~�r�;!��,+��_�����`�v'�˵���C��������NDD��H��N���F����i���Z֨j��=�#�H��М�?x��g:���&�����`nn�p�V�SU��{��]JFty��OM�@�@`����h�M��ǆ��6���0>}���i��u�i~j��o�������	� I�����,}ڪ^��Ou7�%��Q?�,IdY�$ɐe	��@������_��F�VE�Z����h4z�h�(����$���"��:��qqqޥdԯ�� ����(���躎��U��ln�����������s     IDAT�D�	EQ���olwi��F�{##�J�:���ժ88ط��eyG�4�i9DDDto������Q�_k���}�su�$I����n�}uu����R�A����Hľ�u��6M�\�ۛ��������ILN>���٩��sB��.�#z\.7�~|>?�� |>?�~?�͑�L�D��D�VG�z3��V���d3;��H$�����Q����vww���
XZZ�hҿa���XG�Xt ݅��LO��֕J%���~v9o~~��eM���?�%ϑ�zH�e��?���8>~�R�����v�s�V�q(�6�=@�(øݨL"�������m���&�ٌ��.��|��vq�i�X[{�R�[-��sH�:�\��簵�&��&avv>��V�k6����aS�E~�~��w?�^<O����3�l6Q��Q��>|UQ���DGt�E�ӧS�d޾=���	wVz��� �;ln7>4�HFw!
ay��mӥ��x��{���P2��La~~��n}}�BށDD�9���eT����=EQ�2#�`,"""�lp'""z�\.������DD�233�tzز��n���7����n�� Um9���� �4�wz��M��(�x��1���o=�������дv�� �������������I�z���ih4��7Q��P��P��9U��˒�!LMM�zj{�V���6��j��Q?��X\\�$ɶ���css����ӡ�a`u�5*��C�Ȏ���˗��]xr~~���}�Rѯ��޾ Q��m����#R�o����ơHDDD�'��NDD�0I�(�ð��MD4�$I�w�}��z�h6���ֆC���T��s�u�r	���.{�����]|�Q�X���:���P(���Yx���殪*���pw"�	�x���|�x��x<�x��zo~�e�f9<����l��h��l��l��h�Ѩ��l�:у�r�155�D"y�Ǚ�������
�#����n��7P(pr��KK+�D�7t�����Ņ��S�m�כ�&~��/y���ǆ�G�Jq��m�f;�Dźa �b����a�;��(��k����DD��D���b[������+Q���g0<<b[wvv����]z�l
��cՖJ%ll��&��q����8n{�*����`�wy ������|j~�z�p�=p��p��l��S����j��j��j�Ѹib�ijo@Ӵ^G$���G���ӎ�o�T�^���*�J��Q��D"x����v]�in/��>H:=����Ncff֦����*�Ţ#����qz�������Źe�$I������C���������������3MS�u"�n�����Ȩe��i�ᇿd#dE��/
�lkwwwpuu�@*�KO�>���xG��J��l�{���(ff��v�n�!M���͑�2"��(��q��rjz��u�{.(�A���]0�v������_��B�قap�Q��z�����h2�/]\�����,�aaa�h���i66�P.�HFw���.�ۍ�/c����GG��"�����/c�&��7�n�?[#�n�f@͹dDDD�/��NDD�ɲ�i��O�:Q�����/���뵬+�X__s(u��r��o_��nj5M��k�T5�?~���Ɏj+�
66�,ov��%I2�>}����T*����z�ޅdD�4Y��r�4��|�~�k��@��_ҽo�7��A�5h��v[����n���*�m��Ͽ�=]�1�A'������㎚���lboo��P\<��������P���}��Ba,/��>Ǫ������>����X,fYS������0.L �%No�r�\''�,kdY��5M��"Q�a�;��r��TU��u"�n
��XYyA�>������ŅC��7�݊mcZ����ׯ�h4JFw�6M��j��lr�b���go=��0���ǻwoa�f��Q�E�Sû$�?k~E	�(BEH���$CȲ�_^J�i����	�A~o�i�д_NH��=�4��ڇ�:Àa�~�u��㵟}}lhgC��
�1==����^\�����Ω�Y2���܂�u��|{}}�jՁdtW<^��.�˲�4M����Tₗ~2::�gϦ,kL�����U��pz�����F�ٴ*1�^�d��8q*�6�=p�,ok�f�O)� {�����-kt]ǫW߳I�ό��bjjڶ�^�����i�H:h��'���ӎj��:����jY���{LQ<{6���ԭ[�V�����"""H�$�����mo�5���X,t'�T*���َ��UU���*j����H��/�����=8�������S�/_~I�����;�q(}�$�XX���/Q,������,��k���"Q�Q�'��a�z�suS�TD"���\%�"�~?��.LFv*�
<��e�����\;���J�\�a�F���n�����P(�9���2�l�J�p�,w�X�ˍ��(��R����c"""�x��K��;on7M��g���B�Q�^@��c���as��&`aa�pĶ����}G�������,���*vvv p�2�^K��C��1�NN��^ߕ$��8u(�!6�=p�a�E��6M�W`���2M�r��Ö7r=/4MC���}�I��G,����z}E���r��v��x<n[+I2���P*�j�HG���h����( 
uԤ �pS�N��n�V�4w"""�_^�ss��|t��} P�U�������&� ���	<}����V����ר׹(b�<}����m]�R���&�������G,kL�������I�09��(�:���V+���dY��4�O�DDDD}��DDDY���a����AD�M��BD"�S�"�2�4�ӡ��i���J�6u��a���j��P:�+�J��~hr�nVE	CC)T*4�gR�1M�B�B�P�r��_�$	�D�H�J�;Q_E���077��z��/�����agg�V�K	iP����LLLvT�l6������N�ɓ��u�����4Ms u���a~~�v��۷�ܽ��O��Ü���NNN���uE�7u]�w(�)6��XE�OL���:Q7�J%�I�� "�N!g麎b��T*m;'��T*��d3Ǡ�V+P�V�M�"��!4uN|�Z�..Ρ�:��H������`dd���T*q�!�\<���2�ĭ�k��s���ud2 <�y�A���<R�tG��Fkk��0b ��,,�7G����u�C�A�����cYW�V����P*"�"�2&'qz�h48??��E�BӴ?v(�16� @�$�0���9����R)cxx���큮�(�K&#;���^�ch(	��gA�Ǒ�f8�l U�U4�M���=�  �H��l�V�:���U�\B.�E �\��K�  
!�J��n���������4�<yj�s�/i��7o�pp�ϝi�͎Eϟ/"OtT_�װ��j;M��������
$��}cgg�BށTt���l��,NX�{<Q�����u��tvvj;�F����0��DDDD}��DDD 0��E�o����:Q7��
��Ѩe]$E>����>�q�X$b��I��h4���+��D4�C�Z�j�D��&w�0�(��n�qyyUU�Do5IK�e$I�!��%.�!"""G����1,,,"���\���(
]HG�H�e,..۞7T�T����v[�r2�k�$cyy�v�7 ���Ź��6��fg�l�}�ys�\.�P*"��(
&'�z�T�����QK���+E"""�>�w"""�D��a��u"�n+�ˈFc�~A@$���L�[���R����?`Y�(
�� ���JFw��h�\.!�HvԤ�� I{������W��|�z}�z������(��f~Q�D�1<��T*}��y �j������o���z�Ҡq�\XZZA(��b�b����u.�@� `~�9��mm&s���R�mH����(��̡R����}�R�����ץ�ם��`�9�$��a��E"""�>�w"""��0� ��D� ��%�XNZQ��pBR��s�� ���B�e��܂{5�M
$�	H���I8�����M  M�p}}�j��P(Y�;~� �?{w#Gަ���-�}���*Y�Bv� �Ɇ�dA��	`��:h�ņ೯��d�0��ot�� ��<_7Y{��dm�%�}�Ň�����fFd132���/od>@feFF����p8�Tj
�n�zm�I����q��XZZƋ�����a������>�Q�g\.������Z���s88؃�s��$z�j	�dҴ�R)��`�w�����N��aoo�nצTDԋ�(x����BU������}$�bKӴ��_ZDDD��kDDD�s��(뺮o�:Ѱu�]躎H$ҳ�����h�Ѩ۔��0�B�D´i5���Z�ڔ���� ��#�YjP���x<��s6��I�l6p{{�@ ��&�,ˈ���¨�k�t:�JDDD��$I������ڃ&��%���!��c�*��������\.K������>�PSSS��aZ�j�����	�c(O`a��5����E.�'33����ϥ�i�j��ϋ��?�������& ܉���gt]�� �� 8~���J��P(dz8
#�Is��1�i��"��$DQ�Y�DP���j�lJG���v��f�D-M��z�����sl�  ��bJ���,<�nw_ǻ\.LOO��v�R��������$ �Lacc�h�著��Ň���)���/�Alm����Tuu��ӓ!��a	�#X]]7��4��;h��6%#�\.67�L�e
|�xjS*"2�p8�����?��i��8�y�VM����'�DDD�6�џגe�/�n>>���(��H&S��/�<�$	>��L��ddE��E��@"�@��Y�  �!�ϱ!dBi��L&�P(��iZ�v��F���ٌL?Q���jC�v�->���3E�J�(����T(���&��gz���u��4���P.����&[,��Ʀ�����%>}�8�T4,�[[�^o��(�K��~X_߄���Y��v�����Dcdff��o�~]6�A�R�Y#��?�u��)M6��/8����? ����i����_�r��i*6��F�]�Gz։��h4�l6��J�ud���~K�b�8��6��4����B�$�����o���P(�D"�N��F�>ĤDDD4��N'^�Z���+˓�W�V���>������Ҥ������
��h�~G���\]]ڐ����p`{���ϓ�?"���!�k~~�Tʴ����ZՆDDd���ĳg�9��t]���Y��YA����"�܉���TU-ʲ��u]�u"";4�\.�|��u�P�b�vۦddU�R������5�e�P�L���'�a�f��x��z����,#�L�R���nِ�&���(
��s��|p:]}�(
��B�j���ΐ��$�$	ss�X[[7�}�kTUŧOqr�=������"��'1GGGlx�`�$a{�����www8;��q���b� {}��ןmJEDV��>�4l�~)�˚�("���u���)M6�ѯ�e�_k���G����.�R�X��|�F�Ba��ݲ9z
�!�\��T�N'|>�ٌM�h��@.���4oE�D�V�:��u:��ݡ�i#B���\�r�155�ÁZ��"����(A0==���D��L�4p{{���}�Jšd��'�"VV�03cm.��i88�G>�r2A����`0hZ[.�qtt�kVcH�elm��y� �:���˅gϞ�:�D2�=��	�`8�?PU�w<=Ilp'""�_�iZF��?�u=9�,DDv0�JSS�������p���*� �����t�u�p�|�$Y��/��8A@���%�K�Z��7~������c����,˨V�=�^&""��%�acc�d���r P�Tpxx���k�:�ѯ�e��[�F���UU���.�L�����	ӺV����w\p;���W�z�躎��]��A4f�={n:P�~]��G�X�Y#��v:��ƦHDDD4a��NDDD_$I�[]���Q� "�K�Ӂ��#=�|>?�N�7���T*"�HBŞ�?N�6�"��[�X�a�Ö�C�EA�����K���X,"����p����u�(�����p�4��{DDD�W ����?�3]d�k��6>|8Ň�lh��\.�����7��
�o��C�Vr2�����>3�SU;;o�92������M�>~��ADc���bffv�1&����  ��_�4-kS,"""�0lp'""�/�u��,�G�ukc����J��`0��ݳ.� ��@UU���U�n�j�D�ts(F��B�V�)C�\F�QG4�4u;���!�ϱ��~����f��T����p8}/I����t]�g�#��x���_>h���i�������ɔ�����k��?�����y�f�9�d4L��_������=T��,G.�����C
�>|8�)Y577��9��X,�P����e�m����m�DDDD��DDDԓ��8TU��:��J�����(���#�Nۘ��j�Zh�����Fc�T*h�x��5T*�b1���}SR8A>����6$�I�j�p{{�v��@ ��{��Ȳ�h4�h4�f��V�5��DDDd�Ӊ�ŗXZZ���{�cd����s�%YG���E���T*boo�ng��h�B�0���,-�~����~�#A���	��ӳ���`oo�t�1��� ��u��uqqf:H�?�u��M����h������zRU�L�?6#8�,DDv�4�f�D�g��傮�(��6%�~��u��p8ܳN�bq
yt:l�d�V�B�h�,��;�Ο^{��@��jU���@~K�&���t"�J!�^�񳆈�h�H����y���#�}.  �j�����
��sO2�JMamm�h�vn6�����d'�����ֶ�ŵ�>}��͵��!���L�L뎎�����_��(��1�J����+Y��UU��6E"""�	�w"""2�(ʕ�i���s٩�h��t������B(h��6%�~��e8����u�("�!�˲�y�u�]d�Y��a8�SEA<�@�\F�ÿc�2]�Q,����v��v��~�ۍ��i��n�ju~��9I�0;�kk�D�jlo��8==�����H���/`q������NOO�+��s:���~c������>ِ�"byy��o���+\_s�Ѹ	�v�_wyy�n�۳FQ���i�Ȉ���'6��)M�EQ���x���DD�X,"����(��0���`���Ȫb� ������В$#� �IC��ZN2MӐNg��,5!K��d2�f��F�aCB�d�n�L�j>��R���	��|������D�V�W""�1#�"fff����X,ni�򟧪*���p||�ɼd�(�XYY��̬�z�0���)��.����M�elo���6�����ȆT��,ck����z����.L!3� `~~����K�J�L�g�$Ig�n�Ol�DDDD��DDDd�(�E�0�ƨs��0T*e�RS='.ɲ�˅\.kc:�G>�C8����Y�(�Ad2�`�p��#�I�0���N  "��$IB�X�!!M�f����4u����o|
� �ߏ����k�4mHi����
A155�������e:��nqp��b���d��(���B4�T�i�ɤ����MDlll"�� T����qa�[YYC0�Y��:vww��tlJEDVE�1D��QǘX����v{�)��ǚ������&܉����0ފ��'�a���!"zD:�t]G$�Y�����9�oL��|>�X,n:A��r��� ��ٔ��)��C�B!K��`^��|��HdI�Q�����6�`ߍp�mt����B��Fw"""�	��d2���u$��O��f3���G:}]b��    IDAT��9Y��z���>��4��.��vQ*qq�c����X�|aC�����T�;@����Y<{�̴�ÇS
yQ?DQ��-r$�Z�"���Y#�⍪���M����h�񬌈��,�$����_u""�U*�ݞ�u�p�B�ӗƔ��(�H$�'1z�^H��IޏD�TB��F4�Ï�^�O�l4&k�jU����԰n���~����r�Z���GDD4t����7155Y��K��"p}����ԷH$���-8K��f;;oQ�s��c�����Ӧu�n;;��n�lHE�����f�[�P����6�"�~��	�C2藮�.L�(���5M۵)M86��e����(���0ר�٭X,"�L�l��pwww0n=�TUE�\A2�4����*�ՊM�h�j�*�
b�DQ4�w:�H$�(�K\�B�麎b��t��$���=��}zz��'��}c�����gLwy��z����c����dff���Ek�l+�
vwߡ�n9�av���L�t]���5�1Y����������`oo���Ɛ$IXXX�tݐ~�������צHDDD��������"I�����:��t]C��@"��Y�(
�n7�٬Mɨ_�v�z�x´�4���n�V�M�Ǡ�j�X,"�Y�jX�e$I4u4�c�i��<r�,\.�� �FELOOC%��u�:O}A�L�����U��V��'8==E���D� �X^^���s �-������cc�#�L����l�����!w�skk�&U�P�hL�RS������K.//���^�)����֦HDDD������������+��?2�9�,DDvk6��e�@�g���E��E�Z�)���l���"���F�Q68?"�N�\�p�ô^E$	躎J�lCBzL��.2�4��</���O�EQD(��	�^�������O�(bjjkk�H������tpv�	��s,=��(���B,�|���Wx��=�b2�K4��ꚥݞ>|�`:�F�ٳ瘙�5����������_��`nn��]��^�fiz{VӴ�mS$"""z$��NDDD}�$��u��u"�Q(����p�\=���0����c�j�҂A��P���j�lJGä�*��4</<+����x<^
y6�P�Z���nQ����x��1;;�ۃz�U�!-��!I��g����D"	Y��8�n�8::B�R�� =������k��~K��a�ÇS\^^9�%
ccc�(��^]]�s�@ ����M��R	��۔���5;��w�1&����}Y�����������	6�Q�t]�W�(�cNq'���X, �LA����J�Ba��w�u��tԏb� ����׳N��q�E.Zx$�@6���o5d��׋p8�B!�	�� �V��?6�?l�� ��|������E�~�#��o�7�'�خ�]\]]����R����U����^[>T�.�����f�����������zҏ��NNNlHE%�2��^��
��v���MSmJFD�p�\��}���T�Uqwg:�=�i�dS$"""zD��NDDD"I����_u"�Q�4�z�d�g��(�z��dx3z�
y�!ө��("�#�ϱ��)�Jh6��F��nd9�.$I�J\�@w��~�Z������G��z133�?�V��v�=�DDD�DQ<>���u�bqKM��F�4\_���
������LMMcuu��{��lbw���ꐓ�]<��_[ZpS*qxx�E5cnuu�@���������-���ϟϙ^�/�8�����"�#�w"""z]�����?���h�5�MH��`0س���@UUT���Q��@.�C81��'Ib�8r�,T����z��r��h4f��D�e$�)44�c�l6p{{�f���g:��K<����n��n�����h�9�.,,,`uu�p�(>�q4M���%���}5Q�����,O�-
������G��tb{������j{{���sϟ�affƴ���ww�6$"����|��2�[�_gqz{QӴ?�)=2lp'""��$ɩ���3�DD�R*�
�O��#(��9=�CG.�E43m0�e�h�l��ٔ����n!�� �X��-�"�$IB�T�!!=f�z��7h6�_���v��JM!�@�T4��'%""/~���/����@ h�������v6��`8Nlnn#�Y>����Ǉ|>"��`{��n�i����.�s�`++���9�R''�mJED1?����`�����B��?�)=2��GDDDtOE���w�A��F��t��o��Bx���w���nצd�N��_ci[�Z���������H����5D�֛PJ����M!���?����K�����g���rA="��(fg�!
}�#i����k\]]���ݜCԏ`0���K�g����>~�����CNFv�$�ۯ���Mk��6޽��wcg��������4�N����3��O"�p8����QǘX�z��'=kDQ,��)=B��NDDD_EQ��ii�9��FE�4�jU$ɞ��dY���E&��1�K�4
y�����{q8��f30æ�4l�a ��BE�AKǸ\.$	��e޼����j���F�V���1m��EQ�D133�Éz��Fw""�X�;�$������YK�R�D�T\_�����t�ߏ48SS�X[[�,˖�5M����i^/xLDQ��斥ߕ�n;;o��������l�����}��u[RQ�A�������K���W���k�"�#�w"""�*����(��0��#""z�Z��Ͱ��z<h��J�bS2zUUQ*�H$!�b�Z���χl6kS:�K�XD��F$1�v�_ĒL��n�Q��lHHOA�����j�\.���EQD ���,�^/Z�6:������(���������ᗠ��>������<t]`Rz�DQ���2���-�� �w���y���� X[[G$5��4��;l�� ss󘚚6�;;;C:}gC""z�x<�p82��V����g�(�%M���M�����b�;}5EQ<��NDO]�TB0����Y�Q*�n��p�u:T��������ˍ\.gS:�K�VC�TB43���71�bq8�N
�S�l6pww�R�Eq���<�qA������4����.��ƀ�������VWW�D!I���j�p~~���#�E6���9�Nlmm#�Y>�\.cw��<B��+H$��u��coo�&@(����5�B!���S�R�CH������M��8������bm| Qo�(�]�}�BD4J��~��p8zOl����?C�۵)=T4������{�ן��ob>Fn����z���)��8<<��9E ���s�F�'B�i4����32�44M@:""��! �`zz���O�l4���@:��a�G�K�p���P��177������Ghq�%fg��������r�n��z��2==ci��j���{_E���:G��W�w"""I�]���Q� "%M�P�אL&�k=�,��z}�f3���i6h�Z��⦵�@  P.���l��*��n�r���Y[��r��H$Q.���p"#V��F&�F.��$I�z����Eq �aff.��V�DDd;I��J�������Yӝ����u|����'��jJI�KSS�X]]���p?����=...���Fa~~ϟ�Y�4����M A���e���0�����YD�LQ����5./�M�ɲ�Ot]�3�"�#�w"""]��Q��a�Qg!"�V�A
�zֹ�n��R�hS2z�z��n�kiRr(�a(��6$#;��\.�N��H$j�F�,�H&S�t:l����v���r�d2E��EQ�������� TUC��pb""����|��_���*b�x_�M�X��'����u�������啾����6��w��燜�Fav�^X����#noo������WH$�ugg���p�Ѹ{��9<ϨcL�J��L&ݳFż�idS$"""z���NDDD#I����_u"�Q+���S�����M�衪ժ���������Ra��cT�UQ���D-Mi�X���X,0���U�"������n^��$?�������� �2��:t]`b""z�A@4ëWKx�b~�� >��CG.����Ǹ���-:�ۍ����#��)�J���A���Ώ���,^�|e����WW�CND��H$��Ţi]>�Ǉ'6$"����z133;����������[�"�#�}w���h�DQ,�n��GD��)���{�����������P���},.����3K���'���r"�Ӊ������T�U��b��(���x��9�^�W?�����s����*������fff�t~�������WW�h��HHd.�aee�l}1���NOO`\��MMMcii�R���5NO�=	|>޼���{a{���w���i�'�ޫWK�z}��1�J���?��E1��zʦHDDD�p�;�,�u]����s���k�ժH&S=�+E�p����N�b� �����fH4E��E�Z�!�M�4��i8�N�|~K�8�N�R)�ZM4��H�c��nn�Q�V�t:�r��U�A��z�JM!��0�f��&-""�@@8��/����H$�Wc�i��8??�����4MPV�//^,�ի%���t]���1...���F%�����2�̔�d�x����C�W�e�ۯ�(��u�a`oo�;3M�p8�x<9��������Q��i��gS$"""z8�����NŜ���Q� "Ϟ=������ 6�;A����H��W����c��wC�E�355�W��z.f��?��Ǐ0.l!{�|>LO� �LYn��E�4�rY��w(�HHDD����D2�����W-��]�j�ן�ɤ�Ȋl�t:����@ h��v����=.x~�R���W`�v{>����?�&��5�-D"�Z��G4DQ����ދV�ˊ�..�{ֈ�x����=������w"""8Y��������AD4*�2�^/�^o�:��A����_.�E0�Ь# ���l�^�ے��W�UQ*�D!I�.�D"�E��GD���t���N��0x����/���χd2�x<A�l6�	�&b�8_�ի%D"Ȳ�U�ir�,NN�����zm@i���F���چ��|L�T��������(��	���ZZ�\,��>A^�XD*�2�K��pv�ɆDD���$B�ШcL,�0pqqnez�k�vhS,"""z"8������BŌ���Q� "�$�͛oM����p�lֆT��DQ��斥$�a����LƆd4*��7,��vq||�B!?�dD�$�"��fgg��Fڋ����s����Tw"�'��vcjj�dj`�1;���;\__��n�1��!���177�~n�^]]������X,���uK���r{{;�4͆d��b�8��7L�j�޾���{�&�,�X]]�<��~�P����g�$I�������������P(�r�i��u"�q`
�<�ɔ���H$�\.�n�kS:z��I�Orw���q�e�VC�ٰ)!�M�4d2i8��~K�H��d2	EQ�L�2�Fww�(��$��D>Cx�^$������z��!Q�H$���+,.�D0H�P�\���G����X,@Ӹ����tbcc�d
V��5M�����?7�T$���:DQ4��T��>I�^/67�L_�n����w�nG4!fff���Fcb����3��2���w4M;�)=!��NDDDC#Iҍ�iS��AD4.��67�L��޾��t�O�$c{{~���n��qp��|�Ӻ�Tj
�^-Yj|�Q�\���!:���}������4����t:����
�d���8合h�	�BH&����$y ���:2�4��?�V��1�*�bee��X>��h��`�F}��h���666-�ƫ�j��y��:B�e|�����v��3{{�(6%#���r�����U���|>���˞5�$}�4mѦHDDD��p�;��(�4M�G���h\�ZM @(�Y�(
</�ٌ��+��l6�p8b�*��8���ͦM	ij�r�,B�0��c\.R��u�?h44MC�\��ϟQ�U�(�&3� ��� O`vv�����D""�33�X^^���3�|���}I�����%�����d��t���aA�������ڍ �N��`��T�p8������������>1��o 0Z���Gd2i2� �������&}���8?�d:�@��?�u�ܞTDDD��p�"�$Ig��͏:�8Y[�@<7�;;����� Ȳ�����������aoo�Rцd4J�$aii�D��㮮.qv�	�a)�5^���3H&��� �v����4���!Eq �H �L��7?���ǝ=no��� �\�FOQX]]C8�{1���u�>}����!&�q���mi�C�^���[t�]�� ,,����s�u�LGG�6$"�A�x�CſF&����u�Y��UUݴ)=Alp'""���e�/����:�8�$	�|�-<�I����=
y[r��S��o������M�(�K6$�Q������˾���J%���4H=Q��055�W��FwwwH��8���h�DQD8A2�D,� �R����I��j�q��V$���
�ڮK �l6ppp�z�6�d4� ���5�7�������bX_7�ˬ�kx��{h�fC*"�Z� `ee�t�M�2M�ptt`���(���vcS,"""z���NDDDC'�򁪪k��AD4N�n���[�r�i�������f�iS2�Z��_����1��4��;�T*6$�Q��|X[ۀ��|���8==�6�4V</����L��(���0�d2i�ryhZ��DD��A@8F<�@,7�}�]ב��p{{�b�Nk�q"�"�����3�s�4�����cӆ/�|�@���v���f��w���>I<޼�u9��(�Hbzzf�1&����點5�,�UU��M�����b�;��(o������AD4n��666`�Ӭ^�����8)j�8�Nlo���Ȭi���P*mHF�&I��W�'�:.�����	?h���Hd8�~u]G�XD6�A.�c�;� 	��@ �x<�x<����j+���nqww�n�;��&�ǃ��u�|>��躎O�>�����Ѹ���ܲ���n����[�N1A��"��%�2VW�-�A�NUU@׿|R��p,���6F#""�'��DDDdY��?UU�9���������M�r�,�����t���o�r�Lku����~�%=SS�x��DQ�|L�����!*���=����iJ��Ͻ~�ٝ�h��kj������XK&SXZZ�(Zo|�??��[OD0�����=�n�����ln�0kk���ugg�pyyaC""�����DGc�}�|�\.۳F�����������06��-\.�B���h�?��~F���&�Q�Ｑ6y�n7�����t���7��X,ؐ�Ɓ����ں�I�?2����8�aCLG�P"�R���X_�8��u�B�L�B��� ���M�q(�`���\.!��C&��g2�5EQ����h4��q�\��AU���)�#��ذ� ��ncg�-�ͦ�hP�����`o���h`�n��WFc�u:���(��v��5����3"""��,��RUտ<�DD�F���F��� ��ؐ���v���7p8̛�C���r���hH����e�㉾�+��8>>B��R2��'�2����$����_�5��d�
Nv'"�}S{(B,G,��v h4�d�H��8��&B8��ʪ��d?2gg�puu9�d4N"�(��7,-��v;x��-���hP�����M�����;�� �0�^-����:�D��87�"��?WU�o������86����� ��1�1�DD�����7�|I�{�麨RD    IDAT�w�ޢZ������`{�����&�Cӭ`�q��}���}M�V�.NN�#��{�Ɵ��D,G*5�o�7��@�RA6�A.���"zRDQB8F<G4�,��M���"�� ��C�\���(�XXx���g}�j�pxx���OH4�ښ���.vvޢ^�ې�������7���5M�������&L8��;}Y�����Q�A4�0b J��"""����DDDd�V���Q� "G�X���u�N����&������k�M���ظ��x�^�������u\:}���h�6�dD���z�L��L��2Y �:��,�����P���h�EA$E<�@8�k��U���X,"��C.��a��a�x<X]]�{a]6����{�*'7?�x��k���N�����>a'���[8��8�s� фE++kC���T|���J���O�n�?�)܉���vA�a~��#���"�={nZW�U���[�:Z'������kK7U�����H��lHF�BE�x����پ�k�Z8::4�E4NA@$E2�D4Js&p?�,��!�ϡ\.�0��<Ѱy<^�b1D�1�!=��r��t��l�M�4���^�Z�$�����4M�Ǐp{{3�d4n�VV����I��ׯ���������ED555�d25��^�����g� �0� Z��""""�_�!"""���(���u"�qT,������xz�9Nx<d���� t�]�rY�bq�r�^�  ���n�V�ٔ�F�0
��5���M9�,#�J�0�J�2�D��l6��fqss�F�A�r�,5Y%�
� R�)LO����BDt:�:���E�p33�x�r	ss��ÖK��R)����89y���Ϩժ�����(�������U*e���T*1��D"i����ncg�-���hp���#
�V�rY���ڐ����p`nn~������st���5�������o6E""""�	�DDD4A*�a��,�# I޼�^�״�ӥ&������k�\nK���'���r*7���+�D�}W�Vp||���X�,#�!O 	C�3��0�j5�JE��J%Nw'��s�����ÈD�}M��W�QG6�E:}�f�9��!�C<ǫW�P��1�a���+��}�9�355���%X�U�n���󎟓��.�5�{�=4��$M�����ЗU*e|���g�(�u]� �����l�	�DDD4
�,ˊ���������	�y$�Iӆ�P(�f��-�'�����r�Fc�0��(TUE����O��i�d�PU�P��4*�Ӊ��i���M$]�Q�אɤq}��dwn�`'�� �Ӊ`0�d2�����~Ȳ�n��"��(��B����˗�����h^���	�V5u������(�JPUu��CdY����+�x��ׂ�v����}���1����,--�Js{�����[�Z����J&SX\|iZ��t����n׆TD4H~ SSӣ�1�����'���,�S]��ԦXDDDD?�w"""AŢ���Q!"W�`[[�M[t]���[T*ld�4��ۯ��O����O���r*G^����vv�]�J��G�6H��,+���'����}<T�VE�P@�P@�R�dW"�׋p8�H$�`04�F��U�Ր�f��d�j��H$���8��m��fqrr��Oгg���Ţ��F����wh��CNE���iD�� XYY���u�����puuٳFŬ��	�"�܉��hdE�O����8�DD�,�Laeeմ����������p`k������3\\�7�%Q���"fff�:N�5������
 t�qP�h�h�H�8܍*5MC�\B�TB�TD�Vc�;Y�v�
��
��(��>�a(����s��rlj�GG�d,..�=�U�4|����7CJF������w�tx�eҸ\.|�ͷ��k���ɤmHED��L�8��+麎���,�u:�fS,"""��a�;��(�׺��*Q/^,�ٳ�u�Z��}M�lHE��(��ܭ6�_\����lȩh\�b1,-�@Q���+x���a��E�`�h�xGS\B�4T*��JET�5p	���p !#����dI]�Q,�������t���D����
����q�jGG����ZXx����,��j5��3m���#I޼��ҵ �\��`uu}� =vww�����Y#�򩪪K6E""""�6��H9�ο�n���Q� "o��7��L+s�,�&��#�2�����,���\���|��&�Ӊ��U��ᾎSU>�"��R2�Q�����v{ly�n��R��b��R��f�a���xPB����}7�>T���iJ{�X���</�(���/^����a������w_y�_bv����Z����6�O A����h4jZ��fqx�oC*"����B��1�TU��с�Y��-UU�ԦXDDDD��w"""9Y�TU]u"�q&I^��>�ϴ���gg�lHE�&�267�Xkr�d�8>>b��655��ŗ�$���
�<޿�N����q�x<?5����s9��i�\.�\.�R)�V����x<����x�YL �f��J���z� ��W��[k�Z8>>B�\R2g� `yy�d�R}�z�ܮ�ln�D/_��� �Z��ݻ��u�~H4��~?_�:�����
�\�g�,��FUտ`S$"""�_�w"""9�ñ��tv�s"��'���[8�N����C��iRѠI����-˓���<�9��	s��XYYE ��n����d��!%#/��@$A$A8��(�=��i�T*�T����
4M������A������=�����J�
�
�<�ͦm�M4j�(b~~��� �]6����O�>����E	���Ḑy@�\���.��&T*5���ӺN�����6zM���K�p�\��2���6��{.��p8K�v���ш���~�MdDDD4dY��TU����AD4��~?^�~Q�=�Y�u��C�R�)�}��&B����r����=�*o�?U� `v��� �b_��rY������)�8���jx��}7�}�0P��hv�ozo�Z�=?}��(?5������[�V��@��G�P@�\�BFz�� �����z�:��j����bqH�h�ɲ���-�� �˥�۹b�!looCzW뺎w�ޢZ�ؔ��-�Hbzzf�1&���'��mdY�_TU�6E""""�"6�ѸH	�pm��w���&P"����i]���۷߱anB��}�{8l�ɽ^�cww�'�=e�++����}��*���p}}����+I�
��F�D-�2h���Z��R)�Z��Z�p�	ѐI�����������_3� 躆r��|>�|>��wz�DQ�������g�������'��p`ss>��R}�X���M(�ǃ7o��,��b��`�\Ζ\D4x��`ee��{���h�qr�g� �aq \-HDDD#�w"""�,�3UU�p�9��&������M��&޾��nw��h�DQ����Qk۪7����)��q�����?�\.����FcH�&���C8A8A0�}z�Z��O����W�il�#zA���~hd����u����j��R��b��r��`s%Q$ūWKp�\}��tpz��ͫO������k��nK��\GGln�P���͛o-�ޟ>}��ե��hX��,�/;==A�^�Y#I��i�߳)QOlp'""�q�!o���""����D"aZW.�������wg����~��k�y���.�����Խr8���"q� !"8�((w\��.8�MW��KnHD
HAt�A:H����v�g�g��*�d�k���Ņ��ۣk��5���,�{?k��vy�Z���|hۧ$I���FGc����:67?�T*�9�:�ǃ��e���B �����9�������#!�����x��X(�+_��K���"�و~HQx<x<ޯM�^������R�|www����b�PU33����Z>6�����'.�~��n7����ޅ'�J��`��ݫ��,+��x��ߴ6�Jb����]�^/޾��v��w��ӓ'kdY�! xaEDDD=��DDD�St]���z�?�v"�~ �2޽{����t���� ��_�ξ�����Z�0����B�ͩ��I����iLNN�<��T*��� �6�#�O�� �#�� t�ix|�lv��^.�P*����^]w|����x���ۏ?������wwy�j���!�U�Hss�д��]����OH�RmJF����cmm��k���GGG����$I��W������cs������$IX\\����~�eY���C��������g�a���""""j��DDD�k$Y��ͻ5�������������	u ����$fffm՚����m��6��~����������>˲p}}�����٦tD�MQT����C�x<-/(i�(��(��_'��J%��l����i�n7�n�^����(���h �J�򵙝�D��ss�T*���������`��kP�V}"q����6��v�����X�i]�Z�o~�'h4�HED�2:���%��t�WW�O�Ȳ�B4�.��������������'4M��F��v"�~������{�r��GG�MofSo�cnnv>�[����.��t��Qϓeo޼���8Z�%T�T�������	G4@E����@ D ���F.�8�R��Z��\.�T*�Z�p�;�]w��q��t��������r��tu;�W�e�R)����sS�]�i�D�H�$�����͌��/��"�J�)��p8���Ȳ��t���py�hs*j���)�y3Ӵ�4|��oP*�:������p`aa���<�2�4����0���u�������C�����la�;�$EQ�MӜ�v"�~1<<���5c-�����E�#X\\�5!ز,���ɨx�^,,,����|l:}���Oh4mHF4�$I���E @ ������-�B�ZE�\B�\��U�VP�s�%�,M��t��r9�v{�v��r��v�{���0
�(
���C�� !��	Q�<������qc6����wG  ���(m~&������m�Q�D�#XZZnZgY��6��� ������v��wuu�t��߁�����ڡHDDDD�������z����k�?�v"�~��a~~�i���p߁T�.���X^^�:zI�199��ɩ�	��:���p{�jS:���p8����xl5hu�&*�*��
����	��?W*U6���H��������������Ͻ����Y(�+xx(|mh/�� �n#�[�,crr
�����֯=?!��"mz411���Y[�B����F.�f�~���a�����I��@������t;F߫�k��ۅe=�Y��u�]�^��T.""""�z��	�z���S�0�L�s��7of099մ��h�Çߠ\.w �K ����&���K�Z��������P���������}'z�,��������������v�_n��������j�Z��W�^����N�����������p�����ժ(��P���`�F�c�P(��o�?�^kM*����w" ����ξE<>n��0loorq��x<x��;[�=NOOpqqށTD�N��`ii��u;J�;==���ݓ5����a�j�"��?�0ѫ�r�ƫ��eY��?9Q[\\���hӺj����6��9�ǃ����V}&����.�mNF�$���,�����e���
��'0MNp&zI��|nv�mӻ���v�g�,�Z�������Z�F��#=@��]סi����9[���W4�4�?~�0Q{8�y3c��OU�|�t�|>߆dԏdY���"����z�����(�mNF��|�ݟ����~���>}��@*"j�x|���=��b����OO�H�dZ���r����'������z�����a�f�s�I�����Ph�i���>~��e}��ta}}.����B����MNB��u���GZ>�V�������'j'M���������x��z�r��fRv3B44u����~����u4L�h���+'AU��MS�i:4M�������?�YV���T��E�J%�JE<<<�Z�v;���$	ccq�y3Ei�=��'门����5[��j��P�Tڜ��IQT�{�^��im.��������������|��O����ު(�k��ߡHDDDD-�U!�:�$Iw�e�KKDD � �5�u�����xl�W*lm}�C��H$���9h����|GG��>@#��#�2�n�^<���w����4M���0a��������i²�|�`,0���{w(�I���*����?+�$��@�eȲUU��(�/���4�?�4M�Jů��ߋl�%�`0��o�m&��b��O�����Іdԯ�N'��6�v�m՗�%ln~D�Vks2j'n z����uA?��eqqq�d�,�!D  '�Q�b�;�<UU��a��9������������5QUkk����M�������d	�������E,6��B$��8����]׿6�{<^��n���W���m,�c��eY0͟7�?6�7��Ҡ��������K�:=M�r��J��y*��dv.�#�>]�133���і��r�x~~�E��#>�kkk��><��ŝ���⒭��j��������"�v����v��'����N�߇���ǆa�W�EDDD�,lp'""�~ ɲ�B�����x<�{�ݏ��~���I��.��E���B���z�4����\.��dԏ�� ���r�Z>�R���萯-���*<�n\.�n<7�N'x��z�a�T*(��ث�*����2�_�z��X,���Y[�9����>p�����0���!����r9��ns�� x�f��SM��>|��?���iX\\���L� ��y�F��"֡HDDDD��'DDD�t]�������v"�~���ak2�����dRQ;I����E���ت�,GG����js2�G��`rr
���'��i�V��!�EQ�v��r���<6��\.8��g5-=�4MT�T*UT�����_%N�%�~ ss��z�-�h�q||�T��=��FGc��_�$�{��J%qp��EP ���B�:!67?���������� �7��~]�����N����j���C��������DDD�7dY�B4��MDD?322��ť�u�%����|>߁T�n��o055m����GG��D}��vcnn�YM����9./M�Q�e��������������tUz]�Lb�V+�V�_����������x�f����i�����'0�ųQ�k�3l"q���������ʚ��vww�N�;������`ff��1���r�ܓ5����a�s�DDDD�M��NDDD}C���F��mY�a���arr
o��4���ǏQ(p� ��;zi��a�����p�|l�V���	�uI��p8>7�;�p8�p8��88:4M�vLza�a�V��V��V��^C�V���^�eqA� �$	ccqLO�y���b��(
mHG�N�d,.."�.d�������;(J�E���G��Lt u�,�X\\���3�*����i��I���ᘭV�g�IEDDD�m�FDDD}EUտo�_�v"�~577���xӺF���G�\�@*j�Ph++��@>����6�*үRSS����x����p||�b�؆tD�k'��ޝ?��c#��i�u�Y���L�D�^G�QG���ڴ��^��Z�A��Q���B�޾����n�X�0pvv���+.��_�(
��W144d��4M��� �Ͷ9u�����w�ٺ��L�������S��qD"�n��>4���i��m4�C������܉����x%I�Y��u;Q?�$	�˫��Mkk�>|���j�Q��|~���ٞ�T*�����Z��ɨ�y�^�����<�h�T
''4�,�    IDATǨ��/�����$I�4��C��?��}m����UU����o�FB�0�a�04����M����g!8u��~��vcv�-����u|*��=I�X[[���U_�ױ������6'�Np�\x��;[�)��[����B�A�v�17g�I�u�\�O�Ȳ\B�f/�^)Q�QU��0������_ɲ���w���Mk+�
>|�������\.���Z����M�J��OO���[hZ�kM���e�l�$��I�EQ��?�R~�w��@�ȲEQ I���TU�z�ǟ;?I�4MX��0~��4M! ė��i�4۸n���?�������TU���4����j:+��8:��|>߆t4(�^/VW��p8l՗�elm}�"������Ng��B���?p�"I���r��;��{{;h4O֩�����w:�����E��������,�Y!��}k���g4M����V�s�Tć��0�$�vSU��k�M�~��}�l��ɨߩ����7���x�-�J�����ӷ/���~����I^���Iҏk�܀�جn��߱Q��z�$I��͛�g-\�D"����9,���cyy�boQY�P���f��=���bc㽭���J��'���h�D�#�w;�@���F*�|�F��k!�'""����[����/麾o���w;Q�B ��!�BQ��h��:�� ��[N B�ަ�v���x��˲�H$
!
��$�~��}%�����ڞ����i�D��(�h4�suח��?�����~���}������s񺊈zI(���b�X�ψ�$��bkk���X��ѯ��Ǳ��Y��:�d����⢰�(
������5���j���{�*H4`t]���̳v����k��8o��R���4͓�""""z1lp'""��d�恪�U�v"�~e�ryD�#?�D�SN�^�����eY�d2PU~��i�$I���p8��e;���Y�^G2�D�^���o�A��t!���xx(@N�$"""j�ۃ��eLO����-_.����������TA�C�$caa��S������%�(l@H����5�����F?~@�R�@2"ꤩ�i8��w��..�Q�V��QU��4���C�����^܉���oi��GB�� v����4u���#�6mrw��p�\�d2JG���`���`�ש��C0B6�a�15������kȲ����d.I������A�$<<<�������麎��Y,,,��v�||�����	�ـJMi����u���ǜ���촍���$I���2��p�Z!Llmm�X|�@2"�Ph##�ݎ1��w{�$I��p�9�0
�EDDD����NDDD}�4͜������BD��j�J�""�h�T��]�8�{�<<P.�0<�Հ�t:G����h4:�����|��)������,#
at4�4Q*۔�����uP��XYYA li"�T2y���m��ݵ)%�˅��w��|�����mڴG�e~~�VS�e	��(UU133�t�
5gYNOO`Oi�_�����""""zq�vJDDD��#IRβ���P&"��FG���;��Nq~~��L�9�`++kPU�V�a���F>�os2$�P��s-7�Q.�qvv�t����6I�0:������n���y�T*�p:TCCCXZZ��9��h`gg���mNF�433���ɦu�eaoo��������B�n��tWW�'kdY.!� 8������'�Q�k��j!�B����R��F����ᦵ�`�i�P��Z�"�I#��iM�eYF4:�0�����S�Vqss�Z��? Ei�֔�i�D�F�RA�VmSR"""���D������і�� �R)���NO������aii��k�R�`s��E��4H&'�055m���� �T�����+�� ��ƺc ����SX�x�NU��P��:�����-8������,��B�X�s���7�>�#��io �(UU�����D���k~�eYmLF�FUULNNa||����9E�������y3�@ ������9��.!��MTD_H���ٷ���m��簻��0ژ�:mdd��K�jON��H\�9u��(X\\�5P��K$.��f��Q��4ͷ�DDDD�6��NDDDAQ�"����AD4��*���M���(P�T:��:A�����׀��1>�~��l��/d��|�tN�n���s�\.�����r�P(�4�6$%"""�/n�ss�}����3XH�R���B>��BV�MUU���#�}���5��v�Yr���a,--C���ۻ�8���Y�CQW��O���u;�@�Tʸ�L4+�TU�B�d'2�܉��h !���+B��ng!"�|N����I�Gp�Z�ڡt�	�\�zCCöH�\.D"Q��94�$�A�h4p{�B�� �����^�^/���el�"""�W��t���9������>��|;;[����\<H��\.ll���Pڲ,����ɨ�B�VV� ��w�J��8::�@*"��ׇ��n�gg'���O֨�����_w(Q[5BMDDD�?�%IJZ��v;� �$	++knZk>~��b�ɨ�B�!,/�@U��z5�vvvpw�os2D�$!���4t]�9�..�q}ͦ,"""zt]������Q*�prr�\.����5�XYY��X�4�����6��~?���AQ���K�o�����DJ�e,,,��pt;�@�f�H$Ο��e�.����DDD48�����IE�u�i���A��E&�F0l���,ˈD��岜�=`��
��,���l5+Ȳ���(HH����77�0>���&-EQ044���1 @�ȉ�DDD4�4M�������l��S�Z''�8<<@�RnCJt��8���m54@�R�ǏP(ڜ�:���b}}���|>���~V#`���@�c�4qzz!ēu���M!�w(Q�q�;I��b��A�������x��״�Ѩ�Ç(�KHF���VVV�l�J����~Ӈ/D�F�4LLL"�4�F��D"���K����h (����8&'�l��S�a����H�l�,cnn��1�����cgg��������{[��67?�4��Ѡr�ݘ�[x��;����2���5�,'��)�Np'""������i����DD�²2�4���MT*��H$�I�H���4M���u������0���hsBDB�����=����9EA(4���,�B�T�@"""�K��`||++k?k�e	$�7���B>��u=��������ö�������6��������{�޴�T*as�#L����$I��}kk�5W��qy�hZ�(�_B�w Q�p�$$UU��0�ﺝ��h�8�{��Ng��Z���G�Z�@2�x|��omOaj4���A>�os2t>�33�-�$�S�j�H&o��EDDD}��'���m��N�qrr�j�����u	�X^^��� �e�����E��Q7�\.�{���hZ[�V����A�^�@2"���XK�{�ӎ�>�X,>Y����mƟ�L""""��a�;$���V��e�>ʊ��~����l=Ȯժ����<1�������UUmճ��^R(����gMt����DDD��dYA,����f�_���qrrԴ9���Xlss�;�����]d��6'�np:���xokB�Q����J�܁dD�-.���O��r�,..��.I�iYV@�3�����:G�v """�v0�AQ�	˲8ŝ������{D�Q���k�TU��p�t�[��J��\.���a[M�$!���F.�cC1}�j������%�|~�-~��{T$�i�(�KmHJDDD�:I��Ű���H$
Ey�㼇����p~~Ɖ��MdY���"���m7-V�ln~���}��Q7�����ǏP.���h�I����Yh����o�����!���u���u(QGq�$2Y��"�� DD���`}}�V�E�RƇ߳�b@i�������E��lq�?�Y�16����7M6-�J��8G:}�DDD��� ���t�����e���"��}�t�Z�\.����㱿{���vw��h4ژ����p`c�=\.W�Z�0���HFD���add��1���e�k���@# x#����'�� �4M�d���� DD��V�����H�Iax8�L����&R�dYF �u���E�XD�ZisBt�e�P(����F^��YSNu]G$��0�T*�ѝ���:BQ��ű���H$Ei}w�q����c|�t�R���з�������_��\coo��������x��ݴ�4lm}ds;�+�r�199e{�zZ�RA"qѴN���b��Q"u�.���h੪��0�w;� 
�BX]]o��<6�~����X4:���Ȳ��b˲pzzb��]_�&''��ڳ�S��qy�����`s�<M���#��>��xll��8G2y�z�b&&&��͌�fE!�L&ۜ��E�4ll����iZ+����M���u u�$IXXXli1=���bEUU��0��E""""�
6��k�$)aYw�!"j�Ph��k��܋��&w�`����z�XYY���}L&����L�hc2zm~��>�Mc�F��W��L�0�%""�o��:��'��m/�%�Z�D77�B�`Bz�E���"���cj�vv�8�{������w�z}Mk�0������|�Q��bc_wão��f��$ɰ,k@�3�������M^DDD�E	[��;�BD4���
��D"Ѧ��t]G0D:��e�c��u�ަ����rٛ��v�Gpw��z1�e�P����À�緵�EA0D<>]�Q,a���NDDD�s:���~���e�AHR��&�c3���)�Q(�sj;��˅��w���������GT*�6&�nRU�����5on�,�����$#�ns�ܘ�����=�0���4]�����B�a�bu�2���赐dYN!����hP��,/��z�Q(�cs�#�D�$I��������c����.�Y���i��q���CQ�?��4M$�7H$.P��^0!*�ǃ��ID�#�� �h4�H\�����Ņ�a,,,���Q"q���.�`��bcc>��i�cs�6?���$aaaN������9r���CeY�B�u(QWq�;���o��_�v"�AU.�Q.�G�6m8NA�ӷ|>���*�2���mMΖe��4MC>ϭ��e	!pww�d2	I������`&�2�~?���p8�T�0���������~�};��o���z����h�qvv���]����3��/��߾����i�������e��Q7)����u������eagg���D�H,6�`0���T*����(�_B\t Q�q�;�*���c�0~��9��Y$��Ҳ��|>���MNp����-Mtzx(`ww�j����5�u&&&��AQ�e��L&������_,�+	��0��'��L�z��	\__q�+j�Á��[�_T*��l�T*�1u�,?6�����,����.noo;���z�������7�LC�eY���UU���;������x�IDDD�Ͱ$II˲��KDD-�aaa�Vm.����6�����XZZ��p��1�F��{M��%���!G<>U��K�b������Mq�*�+#�2"�(&'��v���\�Z�D777�������X\\��j��������FN�e���#j>����}���$#�^ I��t:�e`�RI��\?Y#�r]�ЙTDDDD��-㩈����QE�u�i��B���b��Z��p�y3�����G&�fC� �,���[!>?$o��^Q���@�4������WI���;\__�^����={���;G022
Y�Q.��x���h�i����I,-�|�v}�j����3�P���#jI�0=����e�׽��x};�dY��� ����J%ۜ��zI<>�@�����z����Ӧ�}�����;�����'p�;�J�,���n� "t��8޾��U{ww���M�&'�����I���e���aoo�z��Ɉ����bjj���e���$�j����&""���r���#�,��t�R��D₻�P�9,-��Ԙh�&����ɤۘ�z��(X]]C0h������ͩ���x<^���w;�@9==�����5�����9ݙDDDDD���DDD�*���g��G��AD�LLLbff�V-��_�ۃ��U�\n����u������ܩ�$IF4����n���_bY2�4./(
/������!`bb
����|�b����s�ӷ/���iCCCX\\ni��r����m���6&�^��*��6���mճ�����eK�<�~�����'��,M��t���M'2�6�ѫ�����{��AD���O`v����B����0M�ͩ��E����ё��K$.pzz����$!ylt�x<�|���<�r� ���������o���z��|�|>���s.ܤ��$	SSӘ��B+��S�� �PU�����5���#��hs*"�5��S��~�H���]���'�4M�{�F���P,"""���w"""z�\�,g��n!"z���`jj�V�����>��h�7����Q��/@�e����屷��!�K
�Ø������J����+$�70.�!""�E�����b�1�����f3��8�.�1��cii	�А�c�899���e�Q�xln��g�����mNED����ޡ�칾���m��Y�KB�! �JDDD���� DDDD]d��z#��׻���5����,��MkB�2�4�HG�T*���
��i��c�NFGGQ,Q�Vۜ��Q�\������i�n�;?B�4!���D�ZC���DDD� bvv��CP��?NB �JbWW���j/�����All�kiׁJ������f3mLF�B�ull���as;�뤪*ff�~���X�RA"���TӴ�n���D""""�I��NDDD������a,u;�k111i{�O�\�Ǐ�sJ�+�(*�DmcY..�qvv�j[6�_�r���#�A���A�����.q{��e��LDD�I�,#�b||����_cR�$�6�S�MLL�͛H��G��L��]��u�����xlճ������~�`0����� �R��UU��a�ӡHDDDD=��DDD��\��j�zjY�OuH�M�P��)�����$I�}L.����CPWh������q8�o>_�^G*��W""�p�\����Š��vzJ�R���%�����	��s8X\\j�Q���#\__�1��Á���p�\�ꏏ�py�hs*"�E������c��ӷ���|�F�$Ӳ�8�TgR�&6qѫgFAQ��eY��Y��^�B��F���Mk5MC8<�L&��W�P( ��!
�n2r�\��\.�R)�9!я	!P(����
�J.���?�|��  ���G�QG�Z}��DDD���P(��o�177�@ �ͻ�<<<�����(
܍�:.cmm��Dn �V����D&�ic2�%N�������æ��D4�4M���[Ȳ���z������׉����B���C�����z'�=�dY�B�����5���0??;O��*>~��j���`�TU���""�HK���\���BpAu���0��'
��6��b��W��Mq��3}�uel,�����,�L�D�HH�:Y�133�x|���2��`F��Q����n�������ɛ��"��43�~���1���1���e�Z�P$"""���w"""��TU��a��n� "zmb���`�#j����^����5���1;��d�6F�\���.��b�5��z16����L=B ������|�:	��##���I� `�&��\^&��
u������JKS�-�qz�    IDAT���	��6&�^�v������i�eY88�G*��@2"�E�H��S����<��N��Y���N���;������ױ������TU������AD��D�#X\\���\������˥$�^�������ҤM!��N�H$ <��/Q��ccc��Ơ�����T*����T
��x�s
�Á��FGc/2� *�
����L�p�5u]<>���ٖQ�jU���Pxzz,�ۍ����>�<6��!�Ju �"�Ӊ���Y�O�L����.���ݨ�����W;�������������ܲ,g�/�䓈�l�D�XZZ��侹����_MӰ�����ᖎ��s���C�^oS2"�$IF8F,6�P(�"��Tw""�G�$!"C8ii�_g!�����52�4,�'��t]���b˟�������0��z�X_MӚ�Z����.2�t�Q/�$	��p�\ݎ2P�d��'kdY.	!� �&�g߾#�`i���B��n!"zm���咭FEQ�D����h��k!����-,K �nXr�\E�\B�RisJ�f,��%�RId�H����M��$I��������	��r��ɲDD�:�\.��O`qq	��8<�77���T*���=\^&����p8���x�^��X����1��!�hc:�5^�����d2O7`�`����c��J%\^&��i����������'��UU��X�v"��(cyy�Լٳ�h`kk�$�^��������D���kA�MɈZ��*"�(��'�v�_謜6KDD�M�e��( P,q}}���L�׌�dY���,���+�����E��Цdԫ� VWנ�j�Z!vv����:���z������\�c˲pp��j��d�����0��C������܉���~���W��s˲��Qcee��Dc�4����|�b_EQ0;���XKǕJ%���T*�)�sI��XCCCx�[w�Z��)�RI�J�>KDD���`dd�舭�M;,K �N���
�������x<,--��?� R�$?q��+4<<��e{�T�0����|>߁dDԫE��⒭Ⱦd���͓5�$5,ˊHw&Q�`��/0�AUUM�/v;�kT�TP(�#�6} +�2��(��
�e6n�&�e!�͢\.#��� t]��h�ir�?��J����noSB��vCQ������#�BQT�6;Q�p8�cqq��������R��q}}���]$�I�j�HK�r��q,/���p�>�0��������B����Wl������ۉ^���)x<�n�(�j����B�?�P,"""���	�DDDDO�e�B1��DD�U ��ں��N˲px�	77�HF���tbii~�����h�۔���Ȳ�h4���1����bY��R�2��`�;�U��D022����\777�f3l ����,,,~��Ǿ��<����X��cnnvZ ����&w� "crr��1��᧦�Gʲ| �X�P$"""���w"""�'躾�h4�,��uQ���M���c$mNE�H�$��O�͛H��_ݍF��H��0�6�ۍ��FGG�i���W�l6�T*�\.�F?""�I�144�H$�H$Y~���k�noS���B�Z}����H$���yh�f�˲pqq���3^˽R�����U�����w4#z�t]����7�G?�N������I�����Z�C�������������4�h4��9��^3����]U�5�_\�����ͩ�W��~,..��r�t\:}���Oh4mJF�2�4���� ������Z��L&�d���ӓƈ��^������(�ё��z��,�\.�T*�L&��_�i��ann�H����*��v9��{�v�����F������'"H���o���x�e���u���B�d��i�M����:�����/�������9Y����=����Ey<��o@���S�$����J)����y����t\�^ǧO�f3mJF���N���18���*�J��ɤ9閈�^���A4E4:����f��nnn�J%�x�����0l��"�J���L�lS2�e�$a~~��1[��z��P*�ڜ���A,6����n�8��Gxxxz�Y�SB� ޸&"""z܉���lp:��r�Z��n� "z�N��7l7�d2���4��C�+�b~~����/��[|�t �0ڔ��I�����^|�;��(�N��J%Q�T^��DD�z8�N��D^��Bd���\#�Ͽ蹉�EUU���"k�8�0px�	���6%�^'�2���ۛ�_�V������D �x�x�v����v�l��E�2KӴ�m4���������V����lRU����n� "z�t]���;�����屽�ŉv�������r�MT�j���c��]�122����n����P����-2�4j�ڋ�������F4E$�}ߊB��d���)^�S_	�������.<��=��v���+�(
VV�
�l՗J%ln~D��kw"z|YXX���ݎ2P���w�^�j��?5���P,"""���w""""���,g�/�%DDD-QUkk����5,?<����F���dԫ$I���4&'�Z�Nuss���#6LQ_�x<���h^[��/ ��E:�f�}��I� P�Րɤ�LޠX,�����I���� o�8˲pqq���3X�զt��TU�|?�o������[ܝ�����~�`��������wO�Ȳ\B��2�lp'"""j����n�^����ADD_&��"�U_.?N,���-`aa	.����*�2���Q(ܷ)Q{I��`0���Q��(�����6�ߢ^�������׵���0d��RI���a��S0����NgKǕ�%������Mɨ8N��o�ޥ)��bwwB�6'#�~�1>>����.���Ӧu��_��j������܉���Z���?2��v;�$cii	�H�V}�Z���T*�6'�^&�2���`bb���puu���c6P_SU�p##�x�[��e����l�L�*�s�������p�p>����oYr�,R������o=�3��RGGG�;J�fn�����p8l��ަ����i�D�������"dY�v��b���`O����?0�/v(�@`�;Q���$�Z�e�i��$I���G,6f��^�ck�#��b��Q��BXXX������R���NO���p8G0:���m˿�Z� ��"����=wA "�g�$���cx8����)­*�KH&�H�����������R���T�U����Mɨ_�|>��m@�4[���W8<<��v"z$�2��Z�ѐ���8C.�{�F�����;��l���9[-.���n�������
�� Ҁ�"��AdRF�Q��h$	&
IP4"!B!
bDDB�������oe�\e������}���v�]�]~�$��}���#]�|��s��B���    P
�   �8ί����[� 𭙙Y��W�Ů�yz��k���mۚ�����HM��0��ζvww�LE{H&�444���A9N�!_�\.��~yy�� <�e)��U�z{��.X֪T*���X��'*
�@3�����)��O�0j{K���v�(�gj�K��ӣ�o��e�U���������܌������1�N>���17���J��[M�  �V(�  <�m������� �oMLLjzz��c��ׇ�:;;kp*<���ZXxU�v����hmmE�|�Aɀ�3C===T�@Ê������Bgge��<�!_ P;ǉ���O}}�J�ze�fC�N�\V&s�L&�|��O�>��������JEkk+:??oP2<'�z��uՏ��:8�op* �MWW�ff�Z�������e��{�q�m�-����&�  h+�  .e�q��o	 x���a-.��jB^���X���A�ᩳm[33��qe���#mnn0am�0�R�Oe�~�vc��a���Rggg��8W�Tj�� ����������_]]]j�[H�JY�LF�̩r����!_h˲5==�t:�Z�2�S������.��eH��477�j���0��ڪ������8�_˶���������ŝǘ�Y��_�usR  �
�   �`Yֿ����� ��������o��rvp����Q��t;%o~~����rYk�
��e����400�����Mv��R��l6�l6���sn�0MK��]���W__�b�Xþ�뺺�8W&���Ź�n����>��/ּ+T�R���*�#���̬��'�:6�O��e�
�s477���d�c��|>����{�s�_s]�lB$  ��D�  ��l����~�� ����I��ۯdYVU�g2��,+�'�s�8-,,���浙̩����ݢxΚYv�@�\N��./����j���v����ק��~uwwW}C�CPj�K�D433��������e��^�z�������}_���l6��d ������:F��}_++����m��z��{�  �-Qp  x��0�0l\� � �d����gU/���޽��r���l��_��ikkSGG�J<�i*�����������y�T��Ņ..�uyy�tw ��m�J�z��{���6Y�V�[Q&�Q&�Q.wI�m?y����u��7(��v���W����x�s��7_+��78�稳3���9��z������ŝ��Q	�pXw   <W�   u`����<��[� ��:::����B���
7�曯U*���E$���+���ռ���\��k|?��0C===���W�@Տ��y���Ź�٬nn��� �3C���/��d���Ŧb����3���)��K�Ԏ��Ŵ���T���Z[[Q�\n@2<G�XL_}�����Q���rI_�;*
N�9�m[������K��紵�y�q������	�   �w  �:�m{��׭� �y�hTo��L���U_�T��7_������𜌌�jff���Ծ����-��^�D"���>���W=��1\�U>�W.w��ˬ��x��b��R�ԗ�Zw�y�B�F�LF��g<��E1Ccc㚚��iZ5�u]W��Lm��$�]z��+E"�������7��7H �I��sJ&�Z��������{w��m�z���7)  @[��  P'�x|�T*m�aXۻ[ ���m[o�|�������}_���uqq��dxN"����400P��|>���U
7H<}�XL�T�������۔��+��r�Ke�Ye�� �-�bquww���[��}�-C�vǌ��3��e(V�EJ$:������`&s���u�n���\���ji�,�����٬�����'�\kdd��1���ζ�ً;�1��aZ�YsR  �7
�   ud����y��� �g��_ipp����0��������M__���j.��a���=moTJ<}��(�J���O������vFx���/.�)hx"����{>Mh�U,k���<O�����uvv&ߧP���4MMLLjbbB�aִ�R�h}}Mgg���s5<<���Ūo�<99���]� ��D�Sss�M������s��ڼ�8�q����u"  �\�  ԙm��<�{�� ��655��ɩ����ۭ�M�,�mkvvN��#5�-n�������$��4�J���ۧT�W�x�i_�P�Q6�U>�S.����I��b�&��������ś�]\����B��%EJ�x�����[x��a���Cmmm����d��U�k���Xo\  ϞeYZ\|�H$��(m��}��,�u�;��m���<�hR,  ���;  @�������  ��622���ꧥkm�ii�y��=ZXXTGGG�k��ϵ��J���X,�iJqJ���M��.};�=�����J�|��} e�:::�������Ӵ	��ma'�����L��g*�JM���S�D533������E�����2ۀdx��vW����w���X���A��x�fff�����migg[��ŝ��Q	�pD��  �&�  �q�?���� ��������%��U���lV�߿��{N���4MMLLjbb�歠=����GP�~�0uuu���_==)%�ɦ~}��u}}�e�{.w)��w ���,K����
�=���m7�F�v����se����)��~}�)3C��iMO�Ȳ�{��Y�������G?W�>˲���V���U���>|x����'��it4��m���R��[��8�w]��5!  ��B�  �Al��G���B�s  ���ե�o���T����͍���w�����٩��W*�^__k}}M�|�ɀ��ŔJ����O�T����c�a���+�r9��9��y~ �S,��t�nut$j��\�U6����m��R�4���Eww����H$j^{}}���]__5 ��H$�����:;;�:�R��ݻ�uu����%	��-4���%�<O++����n����<��7)  ���U.  @����yAu�I @���q}���R<���R��o��Z��M���9z��GI:99���\�m@:�}����n�R����Q2�Ւ7�+����򺺺��'?����D�L&�Lv��3���d�7Q�S����f��f/tuu�.1�l���Ԕ��j}�4|mook��3����N�}�3E�Ѫ�/
���Q�Tjp2 ϝm�Z\|-�qZ�-}���\���cL�,A0$)ߜT   /w  �r�_w]�7[� p?�q���W�������u~~��dx�b���J�j^�y����upp ��P˲������R2٩V��y[z�������n'�{�w��X����Nuv&?�ړ��}�s=��.q�|>�\.�����ݓ&����܃ʁZ__������ۧ��%Y�]���|^��}�͒ �2;;�d���1�������v�=.��˕J�/7!  ��D�  ��l�������V�  ��4----�������0�Ǐ[U�ၗkddT33����Jߕ�崾�����$ڛ�8���QOOJ==)utt�0M�B����+��y]__���ZA�0�j}.�'�]_���xkS��oty����.//)�5J&���_xP1�u]mnn�����.��1��ͩڷ���2��a��C U���p�c��J�����}���l��?<���&�  x�(�  4^�a'a�Z p?�0477���t�k������ʖ��I��hzzF##�5��P�����#�5�"����{�J��J���[�{��onnT(����ձ�-�~��ޡD"��n�};�T**��*����2�r���<�se۶���5:�~����ɱ677����d�5<\}���`_b�. �H&����k��i���X���՝ǘ�y���bsR  �L\�  4A$�W*��_ju @�j��������7p�����/(�HԼ�R�hkk�I�@��b1uw����[]]�J$:�^.�<O��׺������-����� �Ʋluv&�Ht*�H����O˪}Ǖz�P777��s�
헪T(��500���yE"���^__k}}M�|���.����[���T�fkk�]� T�q-.�~�.��_&s����{��D"�R��/M�  ��  �¶��y��ku @���ՒLӬ��b��w�V�Php2<g�ahll\��S�,����lV���Ly�̶�/e���n%�]U?�7Z�*��J﷓���
���0hu<�I3MS��o'�'����T,�t6Y�}_�|�K�=���������Τ�����]}��3���Q���؅;���ꫯ�wTu|ZY��L��� ��ϻN&���ҖJ����Vw?Ƕm��{���7)  ��F�  �y�if� �}d+ �ezzRz��mՓ�<����;e��'�s�D533���귮�V���mnn�u+u��<�������ӣh��b?�T*_J�777*�����Q��c^۶���ёP"�P,S"�P<�!�xZo�T*]]])��T>�S>��*@8����)����8p~~���U��저����iii��]@\�����(�cG  �K��400��h8�    IDATm)C����P�{��i�� $�  �	�֫�   m.��b�\��[� P�x<��o����&��a��͍���zzR��_����<������0������&�'�'W���u]��ܨX,|��~�b��R��Z<[�a~*��Nd���PGGBUߌ�la���ZWWy�r����R�cm�0���555��ǆb����5e�H�v322������	�Ţ���k����z��ݚ��mu��u||����m���<�����	   �  �ζ����?�� ��ض�7oި�'U����C���Q$Ľ���ؘ���e�f��ł>~����@��p�{2��t���~���Oe�����ϋŒJ�b����<�=�+�}�<�)�=ٛJ��2{�X��Օ���t}}�'7����ׯ��9����A���]����s�{����y����^��^hy��<�k`2 �&�ja�,�ju��T(���z�뷖e����M�   =�wZ   ړi���m ψa���S:=V���F-������������lV��뺹�{Ke �c۶:;�J&�J&��L&��Z�j��})���^*�U.���~�#♳m[�h��ؗ�i>��N�X�Tf�)��3�FGG�fg������������XS���7�h�4����X���p� ���r�K�iA��ă8  @Qp  h�q�1���a�\��3��-�߽�Z�[��:}}����P)6C���-��ۀt j�8uu%����gUz�.��U.�T.�U�TT*�T�T��[�\���D"�F��D��F����ߟ���R�����/e���<70O�m;�����h�A;<�JEml������Ў��޾�٧]{���677tp���d ����ԃo�����vu~~v�1�a�㼩T*+M�  �O(T  ��eY������9  �J�ji�lۮ�x�s���{]^f���4-MLLhbbB�aּ��\moo����)��d۶�Nuvv*�H|��9M��)A|*����]�����GE�J�i�πeيD9ND���qE"����y�﫧��}��\���F���_>��<-�aht4���骟�}W�:<<�Ǐ[�.B�R�������:����w�fy @�k�E������ڸ�8۶�c����&D  �Pp  h!˲>��?�� ����;��W_)�~r��ƺ��#��ٹO캹����:�
�Y0��Pz��ޫ�w����?��=ϓ�{��p�N�Ðm������??�?�ؿ��#�|����X,}��~}}�R���` ���ק�ٹ������ٙ��6T,��걓�fJ$����1��<O++�yw�>f����yo�   ?��0  @���R������ /��8z�歺�{�^������M�y��c�<��g�ܤ�<G���'	utt���C�xG[������������"|�}_A|���[�_���|J|?O��mG�q�w�0dY�ÔeY2MS����?U^����bw��	U*�U(T(ܨP(|)�?��� ��ё��ܜR)n�D����ٹ��(g�Y-/�c� �8�^�q�VGi[[[���swc��ᤤ��  �Qp  h1۶���y��� ��3S�z��奖���u+L�vc���G4==�7:�0��񑶷?�R�{x�,�R<���~��P<o�ۍ��|?��������-����0ԧ�Ͽ�~[R��_���O�����W�P�^��X,�P((��O ��rG��SM?�1��\moo������Q�q����R���j}}��5 b����Ht�:J�:;�h���������M�  ���+�   O�m����y���9  ��N�ivv���E�\����tu�op2��v45����:<<��Ύ|���@�1C�X�K��v�{\�X\�h���GU.�U,~.�[b/�J���,���hZ��S���w��|s�Ǐ[r]�	��:;�z��m�;�a��������d �Y:=����V�h[�RIkk+�� k����y��kR,   �
�   OC�i�A�6�g���W�_���4ֻA���5��-j��ѡ��9���=h����a�%���h4�x<�X,���������%U*e�%�JE�E�J����~n�>���yע��iE"��#��jss]777uN��`hhX�U����>|x����'��R��&'�[�m�a���5
w_��Y�`P   -F�  ���D"�R�R��V�  <^"��۷?�zқ�6�x���~���)�?h}�P���Ge2�uN�q�S����{4��{�]�<�S�\V�\V��my�s����Yx�5==����b������x�04==���הJE}��7�&�.�X��kP���C���{\4���r�o4!   �A�  �	�m��{���[� �x���͛����zM.����;U*�&C�2C��iMMM?x��U^[[�����s: ��4ME"QE�E"Q�b1E�QE"�b�O�;����<U*e���JEU*��eU*�OS�)��q�TJ�ӳJ&�Z�y�vww����0�/A$՛7o���]��\.�����uy��,����+E�l��(77���X�w���8�u�_iR,   ܃w   ��4�� �[ �x�ijaᕆ���^S.����;]]����qMNNit4-�x�K?�lV������s: /�i����Ǒ�8�D"r������r�<��~���u]U*�/����~;��B�@���&'�400��3�:99���&%c<Xww����*�T����Hkkk���(�;G̪����Qږ��Z]�p�@˲�}�����   Ow  �'�q�_�<��Ð�(�M���j~~��q��X���Q����uv&577W�.���������Q�r��� ��a_J�x�{�[�-۶d۶l���w[�e�:�����<ϓ�y�}���<��^��R�����S�!b����f444���]y{S�nnn�/����yFu/ņa��������d ^��Ѵ������|T6����0�H$�T.�W�   U��  �E"���R����� ����--��i"��ѡ��י�GI�R���S"����A����@��;�<��� �a��Rxw�o��?LӔm�2C�e�4�O��[����!ٶ#IOb���y
�P��)��w_A(>����/�����o����(�x
l���Ą��1���f;
7���V&sZ�txIL���܂FFF�^㺮�������$ T���G��3������ϵ��s�q�m�{����M�  �Pp  x�l���yޫV�  �O4���ۚ���sz���*&h�����������Dt�u�������_� �|.���_� ��$�C����I����K� Ю,���ظ���|3Q�\�Ǐurr"��v�pyn~uu���ߩ\.50��"�k~~��7{�~�rY��+���e��?�<��4)   j@�  ���3M� ����  O�i���_��p�S����������t:������-��+�]    ?Ͳ,�hbb��ݬ���\��r���`w5 �fY�^)孟F	�Pkk�*wg�f1�aI��$  @-~8�   OG�q�m���H��  �'C����R����WƏ�|�˲444� ��皐�*C��9�0�d2Y���wY��T�W����]__��$b   �l�ijxxDo�|������~a���@�߿��e�kN<��Ȩ���T}�oZ__��ζ�5 @�LO�*�H�:F[;<<P.w���H$�K��݄H   x &�  <q�m�M����V�  �_ww�����49���Dkk+L.D]D�1MNNjxx���g�rY{{�:::��  ��3S��Ú��R$��ɴ�2����6U*��/��Nj��zM�\���;���P?��i�:F[���kss������\���&D  �Qp  x��4O� H�: ��"��޼y�����\]]iy�e�M"��������|�R����1]  ��1C��C���V,{�y�٬��6t}}]�tx���--�Qggg�kr�K-/�W�Ri`2 /Mww���gZ��y����r]���L�<�`Xl�  �Qp  x��=����0�~�6d���g4>>Q�������L洁��ҤR)��̪�3��sPt  x9>�''���|�������ty��c:�t��Z\|%۶�^stt���5�� ��x<���E����(mmkk�ޝ7��#�țr��ڤX   x ��   p� "������ou @cd�Y�J%����0�4M*���"+�J����U(�ٙ��85�öm���k``P��P�i@R   �����A�y�FFFt�(�^nl�kcc��P7�ijvvN��sU�I� ��ڪvv���c۶���e��]��d2�:;��{�m�����k"  ��� 
  ��ض���y_�: �q:;�z��b�X�k�������B��4M���jbbR�H��繹����vUo2  �3488���)utt<�,�rY��;:::dR6�*����7���zM�\����tuu��_ ��a���Wggg����R����UAp�q�m�]��~o�b  ��(�  </ݦiA��=� O��8ZZz���T�k<���ڊ2JĨ/Ӵ�N�5>>��ɜ�t}}���me2gb�  ���0n'�ONN��#���T*�/���Jh@�������Z�mW����R���底&�R��O�����1���+��0M�*�!I��$  �cQp  xf���?[.�������f���g4>>QӺ��}mnn0ugY���G499)�y�D�b����]�}
  ����ib����Olw]W{{�:88P�uL<����ѡ���x^�!�N��:F�������ŝ��Z��<��;M�  �:�  �Y��������� h���a-,,�4����r9}��^�r����RY���Ѵ&&&k���C�RI��{L�  x�>��8>>�h4��󸮫��������:&n�b1--�Q2�U�������L洁� �d�d�fffeTr���\{{;��8���݄H   �#��  �)˲�}ߟlu @�utthi��D�k\����]\�70^�z�]����C�����(=  ���b��Ĥ"�����������5���_�^��m;U�)
Z^~����&�E�Q-,��eU?��+�JZ[[�wh�m�˞�iR,   �w  �g*��K���0� �l��������Դ��`_��l���qG������dY�)��N���ߗ�uL  ��|��K��u�"�v4�a������jy����Xkkk
�q� �h�ei~~Q�X��Q�ZZ__U�X��8�0�a�K�4'   ꉂ;  �3�8ί����[� �<CC�ZXX�iV?*�����*�r��sG��J��d��������������,  @�E"���kt4��I����vvv井:&�/����7���zM��X���Q�x����􌺺�|�����T�ke$�c�J巚	   @�  ���m��<�ku @�ttthi��D�k\���ʲ...��_�=��kgg[�2Ew  �z��b����#��|iwwG�
�v4V*�ҫWK�D"U�)
Z^~����& )����`�c���ˬ��?�{��8�u��	�   � �  �?�4ͣ Z �<�eiaaQ��C5�����Ǐ[
ðAɀ[�hT�yTi*���hww�ޭ�  p�D"���I�0�6���:::���.�v4�a������jy{���D���}�q� @R__���'[���%���(�;�3M�0�1I� 
  ��Qp  h�ht�R�����{I ���Ѵfg�j*_^f����h
�q�N�)��mۏ8S����)���-  �K��ݭ��I���=�<�������h�h4�ׯ_�����5Ah}}M��GL ��N���?��1�/C����X,�y�a^4](�J��y  ���6  @�p��\���V�  4_gg����*�W���<��������ɀoY����QMLLȶ�G����Z��{:==a7  ��`����5>>�d��Q�r]W����ߓ�yuJ�m``@�5=(Z^~����&�[�H����cn�G5��wuvvv�q����뺿لH   h0
�   mĶ���<��: ��,����+ִ���X��klَ��,K��#�P4}Թ*����)Z  |�e��������<g@s�����Y��c5�;;�huu�� �²l-,,>�w-�wy������m�������&D  @Pp  h/�i��A�: �5FFF5??/�0�^S(��ò�����>�0588��ɩ�v�1�����H{{{*�KuJ  ��b1���522��I��RI��{:::TuJ�/�L���75=G�@[[�:8�o`2 ��a���S2�lu��W.����r�p˲�|��ą  @���  �f���b�Ry����, ��xH! C���h{{[Rذl�����!MLL����gu~~���m�����  x�ɤ��1�0����͍��vuzz�0�y�+����lM7l�J%}��� M566����V�h{Ah}}M�b�������B�T��;   �
�   m�q�_s]�7Z� �:�ekqqQ�5����je���r��?�P__�&'��2-����`_gg�Y  ��^;��O�����g������2��:dj�F��ՒzzzjZwvv����<�A� ��it4��/���..��=�q�_u]�7�	   MD�  �Mٶ�۞���V�  ���ظfffj��纮VWWt~~��d�O�����Ĥ��_�*
�����ɱ��]� ��fY���G�N�մc�O���jwwG�l���haaQ��T�&mmm��`��� ��uuuizz��;��~��vv��=ζ��y�m|"   4W�   ��6M�0��V �V"����o�H$jZwrr���5��ߠd�ݒɤ��1=��c��trr���=�J�:%  h�x<���Q����T�q���/����|>W�|@�L���̬�鱚�
}��^���J ?.�i~~Q�e�:J�+��Z[[�wP�eYG��Ib�  @��  �Ƣ��b�Ry�!���Gy �Y,��ؘ��G��Fr�l�RGG�:;�(úd  �?C�T���q���=�l��������r�dR�_/)�i7ah�q���(ǉ�:J�_���*��V1ËF��R�c��  ��(�  �9�q~�u��hu ����?����>�a���mooK��ֱm[CC��P4}���Ţ��utt$�s�  ��>_󌍍+�=�|�JEGG���ߓ�yuH<\:=���Y�Y��u�������&�g�������Q�Έx���me���8�w]��5!   Z��;  �`��o{���Z� �4D"-.�VoooM�٬VV>�R)7(P�0588���	%��9e2����c�  �2��I���jhhH��������������v�A�=�y������r�� ��0MMͨ����Q^�L&����{��m��x��KM�  ���  �2X�iA0��  �����Ą���eտ<ຮVW?�����ـ�uwwk||R}}}u9��Օ�)� ��0S���U*���9�٬�u~δk<���ZXxU�Nb�>~����=���VI��500��/B�P���꽯�|z�k\�r   h{�  ^�X,6S.�W�0�[� �t$�I�~��x���u''�Z__���J�&��T:���аL�|��*��NN�up�ϴH  Pw�HDCC�J���F}��;����P��CB��,����FFFkZW(��ò���� �700�tz��1^�����A�J����pc��L�X�oR4   �w  �$��r�R���� xZL����l�oڕJ%�����2۠d@�"����FGGe��O��)a*�����@���uH  ^.C�TJ������i'������@���!#P�TJ�����jZ��� ����MOϴ:Ƌ���)ݰ�    IDAT�|>w�q�H�*��_iB$   <�  ^�q��뺿�� ����@���5�������AO�eY��hZ�D�.�,�:::����S�   >�F�����b��ʾ?���J��:==Qu9'P�ijjjZ����h�󴾾����ƅ�*ttthnn�.���~��G:>>��8˲�����քH   x"(�  �<�eY���O�: ��F�z�jI===5�+��ZYYQ.Ǆk<=�dR�����2)5C]^^���Pgg�aX��  ������������N� ����ttt�l�]���tuu�իW��;jZwy�������%��D"-,�>�su����潯������&�  �A�  �e�3Ms?��� ��tzL���2�Z�U�:88���&S$�$E"+�S4��9+��NNNtxx�R�X�s ��+�khhX��#u�ި���X���$}��>66^��ajwwG;;��4
��,�����b�x����JEkk+�<���L�,A0*)לd   x*(�  �P�h�����ׄ ���Lv���%�㵽�wss������jP2�q�T�FFF�J��t�P��NN��ɜr�  /�i������tuu���}���P�œ�Ht�ի����i]�T҇����+h=�04;;���d���Ah}}M�b����-�������&E  �B�	  ��D"�y�R�ӭ� x�,���܂���kZ��vv����COZgg�FG��eYu9��y�dNuxx���뺜  <=	�Nkw�.��}_��':88���x�����&&&k��.IGGG��\���J ����Rooo�c���;��8��8۶���y�Q"  �	��  ��ٶ��<���V�  <m��}ZXXT4�i��͵VV>P�œgێFFF4::Z���s������ɜR� �ض���A���*��ߔ�B���������h�D"����5�T*�������A� �v�ozGs��e���w�q�m�m���@"  ����  ��i��At�: �i�m[33��i]������=���0��׫��1���T���|���YF'''����  �3b�z{{544���~��Y��a���s(����9��2�N�533[��A&s���5��۠l P���~��M�:ƋQ(�h}}���DL��A0,�Ҝd   x�(�  @���n���~��y� ��5?� �qjZ��絺�A�B�Aɀ��F���hZ�X�n�T��d2:99���U��  �+�HhhhXCCÊD"u;o�\���T*��v^��b��^�z��ֹ����Ue2�%����������L3x����U*ww���"���r��ڤh   x��R  �$�q��u����9  σ�D���������}�澷�'�	�x.�R=U�@]��.n��dt||D� �' ���@��#����y�0��EV''�:;˰�����Q���ɲ���]\�kuuU�J�A� �a::����ۮ,�[������U��c��U�u�	�   ��Qp  ��m�5����V�  <��Ú���m�5����jmmU�b�AɀƈD"��Ȩ�D�*�����X��'�}���  w�,[���Tooo�of+���H���rݻ'�OM<���+���6���<ml����A� ��b����j~-wxx��ӓ{�s�/���+M�  �g��;   �˰,k����V <�HD����WӺ ������m&X�YJ&���АL��i�w	�@��g:99���9?  4�a�����а��j�L}�Ͽˏ���f�v^�Y���hZ��35�ld�Z]]Q���v O��8��_T$iu�#���Ǐ[�g�� ��	   �w   �Ѐi�;A�[ �<t����k���V�M1�ٶ���a���(�����NOOtzz���뺞 ��(����А�8�-�]]�utt���S��W�s���٩��WJ&�5�_[[[:8�oP2 xӴ4??�x���Q^�R����UAp�q�i�A���kN2   <�  �sl�������ar� �I,���+���jZ�����|�oP:��ɤ���544$�v�z�R����3e2���x� �j%	jppH�x}���<O�̩�Ϛi������Ĥ������VV>�X,6( <�a���U2���(/���Z[�G�0۶�I�u�^��  ����  �e���yޟiu ����i�';e��%�ò,hhhX===���p�BA�̩NOOU(����  �����O��A�b�-��a�l�B''':;��;�x꺻{������ڦA�����ۓ6& ���Ĕz{{[���P[[�U��h����<�כ   �w   �$۶���y��9  �S<���+uw�Լ���X��r]�ɀ�F�������:;;�~�B�F�LF��'*
u??  ���I��5u�Q(����X''ǪT*u??�l�mkffV##�5����Z]���'�'ot4����V�xQtzzr�q�m�5����&D  �3D�   w�,���}��A  ϓa���Ԕìim�R������2J4_"���а����D�~~�� ���ѥ�J��L&���c]__���@�jnn��k� ������]�!S�<m��CM�:Ƌ��]��ǭ{�3���<6���������x<���~��
���P	�@+��RS�4�-"�V���
%BU�.RI�h�T-�BEU�
��a)m�������x<�g�n��>���������<����|?�ו��3���k�A,�[�   �+Pp  ��J��K�^�M��7�  c#�N�O�����Os������T�~ɀx����iU*�*�ʲ,+�sPv �T��̨\.kb"��A�^?S�Z��y�/^�D"���OT.��}��eS�~��:���@����VVV�1V�ݮ��>U_��0�~�+�n�  ��E�   �J$�?~2� ��onn^��.�z��w�vtxx(;ᥱ,[�rY�J��"��_���j���L������"� �a�f�T*�T,���D_j�P�FC�����~�� �V��jssS���� ����;�s��gaj*���u��Q�}O�_�>��0�0�L��^���F   ���  p'�D�O��; ��K$�z���J�{�l^���O�F�+�L�T*kvvN���C9G��S�q�z��TZ ��e����T.ϨT*+�L�<�N['''�VO4�r n�w�������>����ׯ_���! Dob"���W2M3�(c#C��l����ֵ�m���y?2�X   x�(�  ��l��9��~s�9  /��LE����8���ݻ����f�*�gT.�(�J���^��^?����|�i� ��ض�B��R��B� ˲�r�n����S�j�j��C9�����e���޻���y�F���!���R)�z��ОC������m�?�y���    ^ 
�   �۲�=���� xl���������}l�}����j6�CH<-�LF��ff*J��C9Gj6����tvV����  D!�L�P(�X,�P��0�3m���^?S�v��G��\nZ�^}�L&s�ck�Smm���CH ÑH$���7�=H��h�kw�ݭ�L���`UR0�L   x(�  ����	�p8� ��B��W���)��ꉶ��広!$��Q�ݥP�֕�ϯ���Z�!� 0�2�̇R{.��y(�cٶ����]D���������χ� �Ƕmmn~2�����u�mm�V|}g�4�n+�j�I  ����;   �-�J}O����0y>	 ��iZZ]]����~�b<�ӻw;:::T�CJ<=SS9��̨T*+�����nG�z]���j6/n}� �����|~Z�BQ�Bq��^��Z�T��)ha��T*���|���P�����~#���� ��4-mn����D�QƊ�z��Wn�ۇa�eY��y�Ϗ(   ^
I   x۶�c�����s  ^��ɬ��ojrr���^]����Z���CH<e�r�)��3*��J$�Wv�@�fS�ƹ���:���� x�R������Œ���L�ڹ�����jLj�ؚ��ԫW����Խ�m��z��W�
��d���7�����.�y�u����#���7#�  ���;   ̶����>� ���0-..iuu�e�P�jU��on�"�L�r��&�'���������z���Ņ���� 0�,�R>�W�PT>_�v�zR��R;�\�+۶�������{�+C�kggGa��y <?�aheeM���qG;����h�ߺ�q����6�H   x�(�  �1˲�}�_�; �eJ����o>��J�u���V��GCH<�LF��
�����P���t����Z��P� �W*�V�XT�XR.��vI�tڪ���ϘԎ�W��jccC�s��//����O��gmyyE�B1�c�Z=��km�i�J�j�   �BQp  �c�M��� w �KehaaAkkk�,��G_\\�͛�j�)o �tZ�R���8�a�<���t~^W�q�F�!�g�; <g�m+�/�P�~$ɡ�/C]\\�^?S�~�^�7���A&�ѫW�(���E���ig筎��$�ч�YXXT�<w��syy���m����1M�*�I�f   F�   ��8�o�<���0�6 �XK$Z_�P�2{�c�0��ѡvv�R�n8��B��b��B�(˲�z�0uuu�����s5�MA0�s �4-�rS��55�����c�o-��F��~vv&��|�sa��������,ø�Kp�z][[����! ����fg��1vz����>��u5�0|۶��u�_Q4   �P�  	�q���&� ��ozzZ�^}�����<d0���۷�VO��x�L�T>_P�XT�XR"��9���~q�TRx�8����IMO�����d�ÿ��u]���U��u~^�D�[�%�z�J�d���v�]mm�V�q>�d 0Z�RY��Kq�;�����]$�8��w]��G   /w   DƲ��}��Ɲ ���������?h���EC[[���t��x��P.�S�XR�TR*��y}�W�y�F����]]]I��۞ �0e�YMO�5=�Y�]�:����j���ty�?�/J����|�B�x�c��������v�k��P(hyy5�c'Cmo���U�ֵ�e����x�   0(�   R�m���~}�9  �!�Jis��ҽ��@ׅ��_-�J+��+�ϫP(>袒��}_���7��j�n3 p�����ٶ=����f���z�~ƅ��װ,K��+Z\\z�E'gg5�y�F�~o� `�r�i����0����������n]g����<�G	   c�g�   �Z�4�� f� �bQ���(�J����`�w�vt||,&�_�4MMO�U(T(�NO��܃�@�慚ͦ./����R��, |�0��f���45�S.���8#;����y]���j6�
C�H�)�g����d����z]�y��z�>�d �lvJ����cP�������u�iA�,�	   �   `��x�a2�  ��a����W�����)��VK��[j6�CH�L�TJ�|�f�{A�5�)�������+]^6�l^?<����)�,KSSS��?���|���Ņ��3���3=��lvJ���������0utt����ܝ
����d���j��gp�պ�۷۷^Xn�f7�UI�#	  ��A�   C�J�~{����0y�	 �t:���OT(t|�^כ7���Q���0MMM�X,iz:�l6;��a�n���~u�R��i �D"�\.�aB{6;�Q����U���h���)��}%�I����R�}��mm�V�Ӊ8 �+�����+Y�w���������M�X��[<���#�  �1B�   C�8�q]���; `<�%�z�J�d�������C��c"�@�dR�BQ�|A���rg�������͔����[���Se�&'���\N�Db�9��..:??W�q��`0��K`���������`��۷oU��! �+�Jks�l{tw	�5��������k��A�u��b  `Qp  �P9��\���q�  �'˲������e��og�����Cix<C��MO�oӱL��}_�VK��减ܭ�S�N���N)���|��i��g�繺����Ņ��:�<V�<����R��7CjggG��! �+�Ljs�X.�wAh{{�NwC�,�����F   c��;   �ζ��yޯ�; `|MLLhs�����j]�͛7��lF�O�S�'5=�W.7[�]��N�n�uu�R�y=�i� F-�H�ٳ���jjj*�R������T�q��˦.//���l6���W��r:�ټ����;�9J$���$���@��}�F���u�m���y�9�H   c�  0
I�4� (� 0�*����6�L&pt�j���o�j0��6� ����{>_P.��i���Qj�Z��j��j��)�uc��e�m[�LF��Y�r9�rӱ���0��Օ..j4�uq�T��^�D"���uU*�:������m��V#N O��8z����crrr����[י�Y�`I$  `�(�  `$R��Z����0yu +Ӵ�������M�_������UP����,�r9MO�5=����#ޗ2�ݮZ�K�Z-��W������V�DB�̤&''o&�O)�JŚ)C�Z�j4�����e��4������y���ɲ�{����N��!! <�mks�؟'�����{���u�iv� X��W   :
�   ۶������a|�8 ��L&����)�;;oU��D����,K�������t���d��/�E��<��m]]��n����j�(�c�0MLLhb"�a:{6�}H}���Օ./�j6�j6/�y^ܱ��X,is�Ճ˚�z]o޼V�׋8 <-�eis��鉸���N��7o^��w�a�m����/�(   �w   ���8�u��>�  ���崱�J�l�A�7�M�}����f�� |��E����u���L��P�n���Q��R�u��`w4 �m�s%���v�|�r5�j6���l�պ��SS9��o(��=��V����-5��}��,K�41A�=��@[[����d����u���   $Qp  @,��Q��0�  |�R����ƃ'�6moo��nG��]�R��
�9e2=��?����+]]]}(�w��(O�mۚ��hbbB�LF�̤&''�8N��>��s��//����q����ĄVW�T.�<���`�w�vtrr�0� /�u�}S����%�����ku��[�:��]���#�   |�t��  �X�m�g=��θs  �1˲�������NaU�V���[�ˀ8Y��\n�C�=���eYq������N��G�ߋ;0&�RIMLL|(����d&�8��m�<�S�u���~yy)����5�q���������z�@GGG��ّ�s���`����7599w����޾�V�uy�Z۶���A,   �s(�   .�eY۾�� �o�L&����Je�A�����C���2�xBR��M�=��ɬ���/f� ��u�n����n����nw�Y��2S�dR��g��ڟ��/�u���ټ��~u�R�ݑ�dg�)�,K��ZYY}�ϑz��7o����>= ^��r��&'�qG[��{���n]g��� �)��   �  �)�4�� ��;  _fzzZ�<Q�u]������@AD��c����Ie�S�f��f�411�髣��z������Ǯz��z�����_1�l�V*�V:����V*�R:=�T*����H�j��j�.o-��m�!]"�1C��sZ]]S"�;=t:moo���<�t �Qn���ɱNN�o]g�f#�EI��   ��龚  ���H$~���$C;�,  |9C�JE��.���=�����䘢�Ľ/�OM�nJ�YMLL蹼��y�M��Q��������g�0%��/��n������`�f���d�V늻3 �@MJ�    IDAT�<���u���ﺮvw������ ƎaZ[[��T.�(c�⢡w�vn]g� �H�3�~��b   _�y�+  �-�L~�`0�?�0��) �ɲ,KKK�ZZZ�i�ڣ�nkgg[�z=�t �ɶme�YMNf599�Lf��Oz�2a�����}(���}}���ߧ`��X��d2���u���ĞL&���w�����+]]]}(�s��y���Z[�P6����a���P������������v�Jo�l�z��a�eY���Q4   �K=�W�  �bٶ�z��'�� �mR����W477�����h4����Zц02�ahbbBe2MN^O{��� n
���J��zݛ�$1u�c����D"�D��c:�����i���<O�v����R��V��VqG�@�LF++�*�g�G�v�����v�&���0���+����~����O�t���8�����b   _��;   ��q���?w  �"��j}}C����A�xy��2�ɛI�e2��d&d���S�G��r݁\ו������r9�#�I�q%�}~�uB�D�Ԟ|��O�� �n��n_�گ�n_��;��$�I���jvv��w�h4���V��E� ƗaZ^^U>���N�8��ik�S���[�Z��������   nE�   O�m����w  �P(j}}]��䃎�@��G��۽���y?�����0�=�N?�4�\�a����
��=ϕ�y�<��s_L�-�0d۶,˖�|��[��8΋��7u�]u:u���"{[�nGa���K�8	-//k~~���\]]igg[�������ܾ�|�w�������n�o]k��O{��;G   �����3   �#Ӳ�7��� ��3T.�����T*�������1Ew`���T*�LfB��ć���Ąlێ;^�|߿)�{�}�C��Ͻ��s����� ���
�@��+A���P��)�4eY�Ôm[���߷e�_|\���זe���+�u��t>�;��:��z�Ev`L8����E-..ʲ�;���kw��NN���`�����5MOO�e���U�yq�:�4_A�Mq�1   �
�   x��L����W� ϊa������ښ'�=|���ѡ����yn�	<�D�s����T*w�g�����P��Y^�� T�_8�z��}��W�m�S����B�e�z���s�s�����<_/C���E��m�.�o�qeY����������<���ޞ^�EU p�ahuuM�/�����@����L�<�`IRg��   ����  �')�J��_	� w  �˲,---kiiY�i>h�ϊ(�Ӵ�N��N��J��J]L��?���%_�nO�^W�^O�nW�^���(�x/�b{:::һw;<_��۟��Ӫ��o]g�f7�L��v��/   F��;   �,۶�����Ð� �YJ&�ZYY����&��Ew �a��M�������t:�d2���E�S�yއ��K�=Ia�<a�eivvN+++���V����훟;  �r�Sqq�лw;��3÷m�;]����   �w3   �9��{\��	�� ��MLLhuuM��̃�p]WGG���ߗ�Stp�i~���J��L&�L&�H$?|nYV�11�|�S�߿y���n>�}(��!S�ܟiZ��������ۥF���o����*�t ��Qn�������0����0�H���`�G�   xJB   x�l�����X�9  x���)��o<�_�u������%? �2M��P"��P�O$J��7�;�eܗ�y���A_��@�nW�����n�;� ��a�������ڣ��֥޾����E�� �e�.��+���e��z=mm}*��o]k���y�9�X   ���.   �۶���;  Q(��Z]]��D��{}�����䘢;��2M����D�$�8��Q"���׎��0x�%
�P���<}��|}��~���* #e應��d���t:m�{��Z�a: x9(�?��jk�S�[�:��?���o?   �8��   �gö�_�<���� @4����ޥ��kO��G�<I�E��M���x۶eY�l��ÒiZq�+����<��'���y�<�����u���� �1C33���*�J?x�^�����I�0�0! ��ahmm]SS��������^���޺ֶ��y�oA,   ��(�  �9qL��	�`!�   D%�Ή�;���0��
�=>.�[�����dY�LӐeY2MS������R�� P�}_a��|�a(����MYݿ)����Ev����Ny�sg�fgg����T*��}z��޽{���*?�k�����ue�SqGka���7j�Z���m{��oJ�E#   <�  ��L����t�A  ������ʪ������utt(��#L ϛeY��qS�7d��߷,�+���W���<���?�.��(��|�[�%����?.�A� �g; �g��*�Y���*�L>x� ww]n�P6��;����{����[י�Y�`YRg��   �hPp  ���N������A<�� �e�fg�]�q]WGG�:8��Ҳ%   �\Y����9-/�(�H<x�h_����,�����2�ɸ�����C��Vo]g�f'�J��t:G#�   D��;   �%�q���_���c x����VWW�H<�����NN������`aB   `����¢?�9�!\�����v ���r��2�L�Q���iUGG���3�u����/�    )
�   x������g�<� �X�i�R����ڣ�SA�j�D������#L   W"������dYփ����~� �#L /�eY��������5���}w�:�0�D"����_~*    z�   �9��]����s  0l�eivvN��+�*��a���S�����D�   �V*�������e����<W�����ߗ�{&��϶mml�R:��;�ػ�ljg��0�u��8��uݟ~*   `8(�  ��K$b0�P�9  ˲4?����ٶ���B���z�nGWW���   ���d���������og�����C�����(��}ٶ���M�R�������͖� �u�m�?�y�?   0<�  �"8��\���q�  `Tl����Yt���δ���V�2�t   ��e�Y-/��T*�1ocz�����Sl�r��67_)�L�e��z=mm���]H,���|��}#�   w   ��m���y�w  Fɲl-,,hqqQ��x�^�ƹ��vuqqQ:   �v���ZZZQ�Px�>�;�����T |�D"���WJ$�:o0hk�S��{�Z۶���y��b   CG�   /�a����y�7� �����JeV++����vuu���}��V�aD	  ��*�Z^^��T�Q;����PA�G� �S*����+9�w���y�޼y�^�w�Z۶���y�F/�   �E��  ��f�4�� Jq  �ahf����MLL<j��`���#���	  �ǳ,K��sZ\\R*�z�^�^O�:>>R%��NOhccS�m�e�A���-���[ך�y����Ǽ   �w   �D%�4�� ��;  񹞈����l6���|���ɱ��45   �V�DB��ZXX|tq��nk�;@�&&���E�=najgg[�����5M�ySno?   0:�  �"�R���`�O� x�(0  ^�|>���5MM��S�z�\{{���&+   099���%��Td�{k���J{{���N#J ��lvJkk�2M3�(�����F����i��d2�I��=A,   `�(�  ��r��y���a2r  I�\NKK+*��ޫ�l���@gg5�f  �����"{��z�,�d ��MM崺�F������;�0\�q�m0��b   #G�   /�m�����_	ÐW� �199�����3�ޫ�����@���
?�t   x�L�T�<���ee2�G��h4��ݎ./�� |�|>����G�a�8::��i��u�a�e}��ys��   �x�W
   ^�D"�����a�� ��d2---kf���7�]���ɱ4�#J  ���q���iqqQ�D򑻅��ϵ���V�I> ��%---�7j�Sܺ�0��q�e0���   bC�   c������?w  ��t:���%U*��,�Q{A�j�D��t:%  �S411��y�i>��yA�����yd�ۍ(! ����T4?�wܨ�ϴ��w�����!�ulȑ   ��Qp  ��H$j0�Ѹs  �TY����Y---+�|��M��l���@gg5�aAB   ��P>?���%��G�����@��F� �u(�?-��޽۹��&�D��?6�X   @�(�  `�8�����q�  �)3S333ZZZV&�y�~�A_��ǔ�   �1۶U��jqqI�T���u�]���HAD� �u���⒊�R�Qp��j���7w*�[��g}����   �
�   ;�m�U��~G�9  xr����V"�������t||�F�A:   [6���ܼ*��L�z�~�fS��{���"H ��0������|�Qp��nk{{�Nyٶ��<����   �
�   G�m����_w  ��L&���EU*�2M����Z-�Z�*�   *�a�T*inn^���ː�/t���W�uAB �]�����uMMM�7z����^��o=Ķ��<�F   xR(�  `\��i��A|#�   <'�DB����_��8����<U�':8�W�׋ !   *�Hj~~>��z�����D��{���$ ܇eYZ_�P&3w����z��\׽u�mۿ|3�'~2   �i��  �q�0M�MKq �1MS�򌖗W411�����^?�`?   �U.���¢J����o�z=���H��E� p_��h}}S�t:�(��mm��`0�u�eY;��"�_�   K�  0�&M�|A9�   <O��Ţ���#ٱ�����H�����'�  ��,���LE��d2���j�txx��Ӫa� �D"���WJ&�qG�������;ݽ�4�� 6$u��   x�(�   R�f�{.�   <g��T.��4�G����NO�:>>R�Պ !   &''577�JeV�e=z� T��ttt���� #�Nk}}S���7�YnoA�.�b��   ����;    )�N/���_	�`"�,  <w�m�R����R�T${v:m������X��Tw  ���,[333�Tf��Es}�`0P�z������H� <�����6"��	��}_��[�t:��5M�*�W�N��   x�(�   7���7��/�a�}[ ���|~ZK*������3��hD�'  �K��f577���Jde�f��������a${ /�����j$wTC4� �����W��5��H$~u���A4   �ɣ�   |�q����!�o  B�tZss󚛛�mۑ���vu||�j�D�� �=  �;۶U.�haaQ�L&�=}���iU��j�ۑ�	 �N�P��Ҳ�
�S�޾���U�ֵ�a���|�`0�'#�   <�u   |۶������!�q  b�eif�i�*C]\\����I�  `L]�9gnn^�RI�������H� Dkf������c�#ajg�./���5÷,�z��s#�   <�  �/�L&���`��0�~�  I.���¢J�rdS����ժ�����"�  �J$��T����T*�]C5:<<P�~ў ������%�����#ajw��..��5#H$�b����D   �
�   �Wp�����?���  U"�P�2���E%�Ɉv�.fU�'��NAD�  ��0MO���݅���Z=���>
�g����W5==w|���wj4�o]gF�8ο:~r�   �g��   �5L���A��x� �Й��r����MM�"��u�V�:99Q�}پ   ���dT��jvvV���l���KrQ  <�mkmmC�L&�(�������wY:��o���?;   �\Q�   n�8ο��w  ���Ąfg�4;;'�q"۷�i�V����ɤ  ��K$*�gT.�(���@��T�����PWW\  υ�8���T*��;
�������jwY:��]���ag   �3
�   �ض��z���ǝ �qc�J��*�Y
FT/g�j6/U�����*��#�  �qL�T�8��?R�����ժ���? ��i��oFz8�qxx�Z��Nkm���<���C�   <{�  �;J$|0�gq�  `\%�I��T4?��T*پA�^?S�Z��y]aF�7  ����T��jf�"˲"�y0�Z=����nd� F'��juu=������c'wZk���x����M   ��  �{�m���<�ߋ;  ��P>?���y�J�H���j���N�l6#�  ��LLd433�Je6���P�ƅ���tvV�> x�
����V"��ѸO�=�H���`�CC�   ��   ܓeY���+�  @J$�Tf577�t:�ޝN[�ZM''���z��  �W"�P�<�ryF�\.ҽ���NO�:::�� � ��㎁/qrr����;��,������9   �Pp   �q�?��ĝ  |&��jnn^�JE��m�C5���VOtzZ����  Ɓi�*K�TfU("�����3U�U��י� /�aZXXR�T�;
������²��}��9   ��Pp   ȶ��y޿w  �y��R�hnn^�L&ҽ��W�^W�v�z�� "�  ��i�P(�\�Q�X�eEy��n�urr�j�D��F�7  >�ijuuMSS���Ѩ�Nuxxp�����o����C�   �H�  �G�m��=��޸s  �/��dT�̪R�U"��t� �h4T�����dw   �4��T.�U*�dYv��{��Z��j�D�f3ҽ �sGkk����;
��}��m�����C�   �X�  �G�m�g<����s  ��c(��V�2�R��� ��h\�V;U�VSPv `\�������bI�m���Eu����j
�0�� OC*����f�g#�ZM���wZk��Oy��}C�   �h�  �ض��=��mq�   �3MS�bI�ʬ
��#ڗȂ�W�^W�Z�����0�t  ?�0455�ryF339��B5���VOtzz*��"� �LNNjmm=�; gg5ܹ��׸�+   �x�  ��ض�7<���q�   w�L&U*�5;;�������<O���j�ew  ��ϗ�g�8�O��t:��Nurr�^��� ��gz:�����w|�z�L��{wZk����<ﻇ	   �  ���m���y�1�   ��2��*�YU*�C�%����u�a�9  @�>.���3Cz��V��Z=Q�ٌ| ��5;;��ٹ�c�+�����������<�9   06(�   �2l��{��}{�A  ����|��J��R�$Ӵ"?�뺪��tvv�F�\A�dw  �
�4���U,�U*��8N���@ggg:==�����81C��+��qG�W��Nuxxp���m�m��~�#   c��;   =ö�_�<���  ǲ,��e��T4=��aD�rZ�:?o�^��^��u���  ���8*�*�J�����/p�P:=��V������ x�,���ں&''㎂�p�r���<�;�	   ;�  ��0l���������  �hض�b��ryF�Ba(ew)T�u���NO��t:C8  ��T*�|��b�4�����j�S�j�C8 �H&�Z_�P2��;
��}��e����$n�   D��;   0<�m����_w  �єݥ^��z��Z�T�fs(�  `�d2����Ee��!��R; ��2����6d�v�Q��9��z����   w   `�L۶��_w  0��P~��u]���M��    IDATU���h�+��� ���0MMM�\�Q�TV2�ҙ>.��4�t �s4=����Lӌ;
���iUGG�wZk��/���s   `H(�   �g����A�͸�  ��U�=|5��NU���󼡜 ��Ȳ,MO�U.�U,��:)��i���D��U���� _477�Je6���,����y�^��  ����   ��e��?�<���  �F2�T�TV�<�\.7��a���+]\4T����l�\  <U�TZ�bQ�bI��9��&�v:m�j5U�'�v�C; �y3MS�˫����;
�F�z���;���   �w   `t۶��o�;  �d2�ryF�򌦦��z��`���s����h4�y�P� @l�Q>�W�PP�PT"���.//U���V�����\ ���q��mhbb"�(������o^ۧ�   � w   `�۶���y�w  �qT(U.�(���4�7aV
�j]Owo4�uqq�0�x>  �'�ɨP(*�/hzzZ�1����0�Pj?;�����\ ��%�Nkmmc�_�qNN�urr|���e�}���$��   F��;   0z�m����w  /Ӵ���U,U*��8�-@��{Svo���NY �9������ߕ�Dr���}_��NU���󼡞 ��LOOkyyu�2�T���i�m�����v   `�(�   �0l��9��#�   �i0CSSS*K*��J��C?g��V�^g�; �I0C�����ΫX,)��Ұ�����:?��^����\a�| ���\����b�1p���}�j�;��m��o��    F��;   ö��<�7�  <=���*��*K�����<�S�����������  LLLhz:�aR�m�C?g�}���3��gj�ZC? �e3CKK+*
qG�-��vu~^��Z۶���y�}ȑ    |
�   @�۶�o��~K�A  �ӕL�T(T,�T(�eÿݽ�tqq�F���˦�����	 x���r�����
���������.//U�_�ڹ� �v����L&w|�0����F��N�m��k��}�c   ��  �'��s�� ���ޝG[��}���>��Sթ�n�����2
Q�AA��2�t�4�(+D�2&*�S��jE�!�6ѥ(D����j�]�tk�3���)Tݺ�����SU��g�|��k�S�<�|Ww���}�o?x_y����r,/��ť=9�6"bgg����=��p�'?���כ����X\|rJ{�?�����?��������(�rO~. G���d������u��/������/s  �>� �>��#O��� ��H�$fffbaa1������\��-����x��Q�����Ǐb00�@DQ177��󱰰���{����6�������x�x5ڶٳ��Ѳ���Ͽi:�O��ŵmW�\����#�����WU�[Ɯ  ���;  �#y��PUU_�u p0E���������M���~k����aTU�g?��dYsss����t�}&��姲,�~�ȣx���7[�'N�:'N��:���4M\�r9��VGZ�����7  ��w  �g�����,{� �A����l,--���R���E������mcss3VW���j���:8$&&&���>??��3{��/�������x��A���G۶{� M�x��b~~���G�4q���X__i}Q*��?s  �� `ʲ��u��]w  �G�e����d���嘘ػ��#"��a���?z_[[3�p ���φ����cjjzO�;Oi��~��=�� ��^�������]��>꺎K�>���#�ϲ�{���1g  �d�  ��,�������; ��iff&���cqq)������ݷ�u��k�Nx___�������eY��s1??�����Ȳ|Oڶ����x��a<|�066F;y �evv..\x=�,�:��QUe\������i}Q�]��s  �� �>�����p8�#]w  �[�f1??��K177sss{>�޶mloo�����������������=7�>;;i��y���v<z����aTU�� �^����ٳ�������q���c0��>��着ꏎ9  xA��  `����;���c]w  GG�籰�������ӝt���<;�}}}=66֣i�NZ �4Mcff&fg�bvv6���ߟ�ekk3=z�?�ǏGU��t ����i�={.����Na�� .^�x�Ñ��y�G����1g  /��;   y��᪪��; ���(�XXX|��.�u���������uC� �,I�������٘��}�����ONT]]}�=���|�* t�(�x��7bj��7��;;;;q��ǣ,Gz�\[�,����  ��  p@E���7�� t������B,..���R����Z�z_]]������X��ͭ�h;k�k��ĳSٟ�i&�4���=�����Z `7��g�ף(��S���V\�􉨪�}�&IҦi�{���=H  ^��  8@���֪���m[�� ����d,,,���b��/D��봧��g����������J�И��������\���F��6�5�������N{ �E,/��g�E���zlnnĥK����]�$I[�>?�i  �+��  �^��MeY���m��ly ����O������������[�eY���Zlll���flnn���V���ށ�)I�������阙�y����MD�������3��Vc{{��$ xai��ٳ�cii��F���W�\��i�wm�$uQ�u8�_{�  �"� � ��������m��1}  #Ȳ,���b~~!���c~~.�4�:+ڶ�����܌���g'��îӀ#&�󘞞�����1;;�o�]����l����GQ�e�Y �JE��������:�=z�(�]�2қ��$��,����~b�  �WȀ;  PEQ|~UU?ٶm��� �B�$155�t�}>bb��u�3UU���fll�?~ߌ����N��$I�������٘�������'�N{�,����뱺�8VWW���Ciff&.\x=��:�ݿ/nܸ>��$I�y�qY��  �10�  X�����,�e۶�g" �LNN>x������鮓�ӶMlnn����������ފ����Ӏ}jb�SSSOOd���陘���$I�N{���V�������X]]���� `얗��ٳ�"I�Lw�މ[�n��6Mӭ<�?g8~l�Y  ���Z ����1�M�4�]�  �*y^���l�������^o�}pM]ױ��[[�?����xG@��199SS�155��199Y�u��.��0���c}}��sY�]g��I�4Ν{-�Nan޼���im���^�vvv��9  #�  p8�H���M�,w 0.����a�٘������(���Oi8���f��l���flmm���N��lw��R���٧��������tLNN�ۓ_뺎�����X������X���ͮ� �3���oD�?�u
#j�6�_�>i}��������m  ط��]W  �Ȩi���iNv �W&''�q������xj�;�e��I�[[[������N}��i��dLN�crr�'�O��7�DD4M���8�}=������}c~~>Ο���x[۶q���X]}<��4Mo6M�K#b}�e  �^0�  ��d�e�����C  ��$ILMM����ﳳ���i�i#��*���cgg;vvv�}�����N�m�u"ho����OF�����d?��~��Mڶ���g��뱶�m�2 �ɒ$�S�N��ʉ�S؅�i��勱�>ڬz�����"b0�2  `���;�  �n�y�����  G^��1==33�1==��3133��Od�dM�����'��<;�����sY��c`��!�~�`���,css#666bss367�<�� xy��k�����]��u]�ŋckks��y��몪>7"��  ��w  8��<����/�: `���z13������tLMMG��ۦeY���v�vb0�p8���퇡X�4Mcbb"z�����<OL�����Q��3_H۶�����a���!� �"��g��ܛZ���p/~|�߁�<�����l�Y  @�+5  �H�����,��� ��"I�������駧�����T���]��M��p8���1c{{;����a�'ϰ��4}:��{:��:�ދ~���E��5��������X������ڌ��uo@�Wdy�X�={���q����َ�?eY���(��S��7�9  �+:  8��<����;  �^�����০�"���^������>�,�(���������m���)����zQ��G��{�޳Sس,�:����*�����̾��d���]�����Y�?>�Na�66����KQ��H����c�  :d�  ��<Ͽ����� ���z155��S��������D۶Oއ1��4 ��@|YVQוS��4M#��C��=�����[wTNM���y6���c� ; �~�.�qd~?LVW�իWF�Nxz����9  ��Ѹ�  DQ�����ض��  �1K�4��&cjj:��~LOO?~?�'U�V�4QUUTՓ����~�\E]��X��ߕeeYF��߭4M#ϋ(�'C�y^D��O�<��(�����{�go�;��V�m��`���O�׷��ck�ɩ죞4
 ����R�={>�4�:�]��^ܸq}��I�4y���,��x�  ���`  !�^�˲���mMU t"�~�ٰ���dLNNF�?�~�Ȝx��ڶ��n�i��?������m#����6����m�̿����m�>[���Z����S�}2��dh�ݿn�y��_o���e��z2L�D�$�eٳA���β,�$y6t��E$ID�呦����^�_۶���;;۱����4������y�� `�H�4Μ9��ǺN�����x���#�M����z_3><�,  `��j	  1y�a�4��i�^�-  </������zr���d�yp�UU���φ���z{{'C� pPLLLąo��ߑ��m�ƍ�������'I2���Kʲ��1�  ��w  8�z�ާWU������ �Ѥi��ĳa�'��O�����,�!=жM����y:����T�����<� 8X��������{ 5MW�\���Ց֧i�Y���_s  ��p �#jjj����οo�f��  ^^�7�?z����'��]��]g�k�'���� ���� vv�< �S�$q���8~|��^@]Wq�ҥ���i}������̈�3�2  `?2�  G�B��m��t�!  ��;O���&������䳯������j�������������?��ى���T ��^/^{��������p8�K�>������eٕ��?3"6�[  �W� �<�󟩪곻 �{Y����DE/z�"��EQD������(�"�f�S)�a�eeY�pX>�~8|�χ1�1�D]�]� ����B�?�ZdY�u
/`kk+.]�UU��>�󟯪�s"�o  ��y�  ��H�<�UU}E�!  $�s���5����E�yY�G��]G�꺊����������Z~��i� ��H�4N�:Ǐ�t��Z__�˗/Gӌ�f�,�>\��os  p p  �ɲ���u����  �p����㭡���Ϟ����dY���]��:���p��A��o���߿{ �^���ǅ����d�)������עmG{���{�s  p@p  ����_U�w��  ��4M�>�H�4�,}��G��ӓ���<�$�,{k]���i�~�?7{ן%ID�����'������iڨ�w�TY�U|�O�4�:ղi�h����5Q����m��?yn�'�ܷ~f۾��i��� `YZZ��gϿ�w2�7߼o�y{��I��Y�������1g  ��  �]z��7�e�7ڶ�*    0vi�ƹs�cqq��^P۶q���x���H�$i�����p��ǜ  0� �������u�۶-�n    �~�.��~��^P��q���X__i}�$�,�~}UU�l�i  �d�  ��z�ާWU������    8|�������>L�*�2.]�Dloo��>Mӵ�(>{0\s  p@p  �ϱ4M�]�4'�    �<��ܹ�1?��u
/a{{;.]�D�e9��4Mo7M��p�e  �Af�  �T�e����O�:    8�fff��.DQ]������ʕ�Q��H��<����~eD�[  t� �Q%y������u    p�$I'N��'NF�W8�<�7n\��mGZ�e�G���1g  �D�u   pp4M�,�Vڶ��]�     G�׋7��@,--n?��|�vܺus��EQ�骪�e�I  �!c�  ؕ�m?R��m�<|*    �>�7>-&&�]�����+W.Ń�GZ�$I[��/��Ɯ  2�Q  �211����Gڶͻn    ��4����s����u
/�,˸|�blmm��>I����}�`0��1�  ��w  ���z�Ϩ��g����    �?�����^�����SxI;;�q����#�O�t#�����a�i  �!e�  xY'�4���iV�    ��$I�����'OE�I8�����ʕ��4�H��4��4�/����-  3W�  ��0�������u    t������bff��^��Ǎףmۑ��y����1�Q�   ��w  �UI�<�HUU���    `o---�ٳg#M��SxIm�ƭ[7�޽�#�ɲ��u]��1f  G�+K  ��i��CY�k���n    �/˲8�B�<y2�$�:���4M\�r9=z8�6��?Q�����  8Z��  �rEQ|sUU�׶�W�    ��������/DQ]��
�e�.]����'I��y��ʲ�cN  ��  �X�y�����GM���n    ^�4M���S��r��^���͸|�RTU9��4M��,��eY���  �#Ȁ;  06���g���n��X�-    ����'��.���d�)�"�=��ׯF�4#�O��N�4�<"�o  pTp  �m"�󟩪�?�:    x1I���ʉ8y�T$�Q�����[q���s�y��۪�>/"��  �:W�  ��(��o�e�;��     v������bff��^��i���+���x�=EQ�@Y��}�Y   �u   M��`��Y�4�&��    ���c�������SxEʲ�K�>�#�O�����;����cN  �C%  ���z��,��o��n   `�*�^�?>fg�N���ڌ˗/EY�#�O��*������9  ��  ��+����gM�Lu�    <oaa1Ν;Y�w��+��ѣ�~�j4M3��4M��<���p��1�  <ǀ;  Е�4M�i��]�     y�ǹs�c~~��^��m���[q��dYv���ώ���  �7�  @��<�?RU�o�:    �����8w�(���^������+��6��z��?QU՗G�hG�  �bY�  ���4͇z��d]�_�u    5Y�Źs����g"ˌ&;;;q���ckks�-m�����o��v�i   �('�  �B�����,�϶m��    {������Z\�z9�i}�$UQ�8�Θ�   ޗw  `���z�UU�O5M3�u    VY����gby�X�)���{w�֭�Ѷ���z��_8?:�4  ��p  ���,�~���7�   ��fnn>Ν;���C�i��q�Z<|�p�=Y�]����#bu|e   �c�  ؏�,��^]�_�u    Y��ٳgcqq��Ơ,�q�����yO�e����/��юz  �#Y�   �mۿ���zu]qxs.    �������>-��g�Na677���O�`0i}�$m���Y����9  ��  ��^��eY~�mۼ�    8H��~�ݻw7nݺm;�!�I���^�����ǜ  ���  �����/)��_4M��u    ss�q���(���Ơi��q�z<|�`�=i�>,�����b=Kg    IDAT'Ƙ  ���  E?�󟮪�Wt    �U�q��XXX�:�1)�2._�[[�#�����TU�1_  ��a�  8P�,��u]{�    ��,,,�ٳ�"��S�����r�rTU9�,��B]׿o�Y   ��w  ��)��wUU��m�f]�    @�z�^�;w>fg�Na�<�7n\��mGZ�$IUŷ�ÿ9�4  �Wʀ;  p �z�Ϫ��7M�U;    ����cq�̙HSgAVM�č����#�I�t-��/��n�i   ca�  8�f�<�UU}F�!    ����~�;�ZLOOw���ø|�bloo��'M�_h��s#bc|e   �c�  8蒢(�VY����    �$Ibe�D�<y*��K�����Z\�v%��yOQ?�^)  pй�  �<��P]��m۴�    ����8w�|���]�0fw�މ[�n��>I�:M��[����1  `Op  ��(>����4�L�-    �dY'O��cǎ;�����*�]�kkk#�I�t#˲��,�5�4  �=��  8lf�<�骪>��    xYss�q�ܹ(�^�)����V\�|)����{�<�hUU_�+  �[� �C�(��)��ۺ�    �QE�9s6�Na<|�0nܸMӌ�'˲���[ǘ  �	�  ��U�QU���m�u�    �Z^>�O��,s[�k�&n޼�yO�$UQ�2���   :c�  8�z�ާWU��M�8�
   �}�ߟ�s�����t�)��p�/_�����i��(�/���   :e�  8
�y��DUU_�u    |�4M���Sq��J$��񏂵�ոz�J�u=�<���=����   ����  ���j��E1�4��7�   �O����o|Z���n?ڶ�;wތ�ׯE۶#o��z�kY�_�O�  P�� �#���}MY�?жm�u    GWQq�ԙXZZ�:�=RUU\�z9���Gޓ$ɠ��}�`0��1�  �+� ���L��?�4͙�C    8Z�$�cǎǩS�"M}��Q���W�^��,Gޓ��~���[[[�Ƙ  ��p  ��$��[U��u   ��055gϞ�����S�Cw�މ۷oE۶#�ɲ���u�5ь�  `2�  iEQ��UU���m�   �XdY'O����W�NaUU׮]������$IR�i�_�u��ǘ  ��p  ��^��YUU�d�4]�    p�,/�S�NG��]���677�ʕ�Q���{�4}P��_c  ��g�  ��"��XU՗t   ��755gΜ����S�c��ݍ[�nF۶#���������1_  ���u   �O4M���<ϋ�muxC0    / ��8{�\�={>z�^�9졺�����q�޽��$I��y�?VU��Q��  ��0�  �I�<���i>�4�T�-    I����r�:u:�<�:�=���W�\��p0�4M7�4�UU�?cL  8p�  ���4M�i�_�u    ����L�={.��ɮS���{w�֭�Ѷ��{�<�XUU_��+  8��  �"�,��u]{�    �?EQĩSgbii��:PUU\�v%���Fޓ$I����-���1  �@3�  �>&&&�r8�ݶm�]�    н$I�ر�q�ԩHӬ�:���W�^��,Gޓ��NQ_;~l�i   �w  ��K������%]�    Н���8s�\���B8�ڶ�;wތ;wތ�mGޗ��Ǫ��x<�:  ����;  �.E��eY~0\O   )q��٘���:���eW�\��͍�lk�,��u]p\]   ���  �]����M���۶uL   �!��i��������i�9tdmm5�]�UU��'Mӝ�(�v0���   �   /�X��?�4�/�:   ��XXX�3g�FQ]�Б�m�֭�q���]����cUU}aD<O  ��e�  �%E��eY~0\_   �8{�l���u�B�vvv���+�����mm�e�����  �3�  �&&&~�p8���m�]�    ��,��'OƱc�#I��~�=xp?n޼Mӌ�'Mӝ�(�v0���   =W�   ��r����i���:   ��I�$����ԩӑ�y�9t���q�Z<z�hW��<�hUU_��)  8:��   ��m�b�כn��W�7   ������o���HӴ�:���/~<677Gޓ$I����TY�_���  .   ^�<�U�4?�4�\�-    ��~��O������S�X۶q�Λq�ΛѶ����4]˲��˲�c�  8r�  �G?������t   ���<�'NƱc�#I�d~��øz�Jlnn�j_��?SU՗F��X�   �0W�   cT����3m�f]�    eI�ıc����S�en����~�Z�u=�$I�<��pY�f�i   G�w  �1�����ʲ�ɦiNv�   p-,,���g���u��>P�uܸq==z��}i��)��K��/�)  �0�  �W��(�FY���u   �Q1==�O���陮S�'677�ڵ+1v�/˲�u��ь�  ��p  �CEQ|sUU�۶m�u   �a511�N����ŮS�'ڶ�;wތ;wތ�mGޗ$ɠ(��9x�y   ��w  ��w"M��4��u   �a��y������W"I��;;;q������վ<�?VU�Gă�  �^��   ��Ͷm�\��+������c   ����i?�.������y����q�ʥ(���{�$i{�ޟ*��k"b{|u   �W�   *��s�����Y�   � ZXX�ӧ�D���:�}��ʸv�Z����j_���,���,nLi   ��   �+�,�������   ��bnn>N�:���]���<~�8nܸUU�j_��?VU�WED=�2   Fa�  `���z�����k�f��   ��jzz&N�>��3]����u7oވ��j_�$��(�e8��1�  ��  ���<��qUU��u   �~������S����u
����F\�v5�����y�����("��  ��ʺ   �9�M���<ϳ�muxc2   p��z�8}�L�;w>&''��a�i�&n߾ׯ_���Gޗ$I������F���
  �-�   �TQ�[���7M��u   �^��<VVN���+�$^��ݶ�6�ڵ������}i���������0�4   ^��    �[Z�_/��   �Y�����cee%�ԇ��nm�ƽ{w���[Ѷ���y�CUU}}D4�  �ep  8 &&&��,�l�f��   �qH�4�;'N��,3��{��ىk׮���֮��i����o����ǔ  �+b�  �������UU��   xU�$����8y�TE�u�؃�����4�;|=�󟪪��G��x�   x��  0Y�}[�4�m[��   ���R�<y:z�^�)�c�� �^����ڗ$�0���[��_S   c`�  �`:����UU�˻   ح���8}�lLNNv��>������_�S  ��p  8��<������m۬�   ��3==�N������S���a\�v566�w�/I�:˲?ZU՟S   cf�  ��������,�Q�4�n   x/SS�q�ԩ����:����{q���]�ڞ��͢(�t0|bLi   ��   �C�e���4ͷ�m�Z   �&''�ĉ�����u
�K����y�g˲�oǔ  �2�   p�E�9u]�h�4ǻn   ��~2N�4���<�7o�x�S���y����Ϗ)  �=f�  ��I�,�KM�|���  ��������S�ً��m�e�W���ED;�4   :b�  ��*�����H�4�]�    �[�ߏ������I�ehF���?Ȳ�7�e�/ǔ  @��Y   8��,��J]׿��   ��1�΋q���:�=������#bwS�   �0   y�I�4?�4�B�-   ��g��Ѷmܿ/n߾�"��?N�������1�  �O��   pty�UU_�u   p0�����r�`;����׮]����]�����������_}   ��;   G����W�e��M��t�   ���q���XXX�:��m۸w�nܾ}+ڶ���4MW�4�������   ؇�  MNs   ޗ�v^���f\�~5vvvv�7˲�u�[#b���   ���  ay��ڦi~�i���[   ��czz&N�8ss�]�p 5Mo�y;�ݻ�"��?zzj�?O   ��w   �,˾���o	׉   p����ŉ'bff�������~�Z��>x�����������ǐ  �ap  ���(�����M��   �;I����B�8q"&'���ဪ�*nݺ>���4M�i��UU��1�  p�p  ���,��R�4�޶�kF   8Ē$����XY9�~���Ǐōף���nm�,��u]sD4cH  � 2�   ��E�u]���iV�n   ^�4�byy9VVNDQ]�p��ø~�Z����zo�eo�i�eY��1�  p�p  �SI�,���i��i�   p��yǎ���W"˲�s8�ڶ������۷�ivw�z�$M�e�[UUpLy   p   �E�z�O���G뺾�u�OQ��EdYI�D۶�4u�eUUE۶]g  h��D�������HӴ������~�jloo�zo��7�<���p��ǐ  �!a�  ���y����ڶu���$ILMM���LLNN���T�z�H�_��D۶Q�eloo���vlll��憡w  �LNN����XXXx��/x?MS��۷���{��.O��β����;�S  �a�.   �q*��TU�˻a�K�4���caa1fg�^�)�M����F<~�(VWG]ׯ�  pX������ɘ���:�Cbmm5�_�e9���<�?ZU՗E��W_  �ad�  �]+��[����m���na����q��J,..����O�i�x��qܻw7������   �����XY9���]�pH�e7n\���ǻޛ$� ��?P��_C   ��w   ^�l��?\Uկ�:��arr2N�:ss����͍�{����  pP%I��K��r"�}�C��h�6�߿�oߎ���'��y�O���ʈ�|�u   v�  x)_U�凚���GTQq���X\\�:%""�Aܻw7>|M�t�  0i����r���DQ������܌7��������i�V�7��!  �#;   �BQ��UU��mۺ�<B�;�N��,˺Ny������{q�������  �W���űc�cy�ؾ����:n߾�������O��������   ��   xe�<�¦i~�i��]�0^y�������|�)�m�x��Qܽ�f���t�  �B&'����X\\�$�2/���Ǐ�ƍ/��4MofY�[ʲ��1�  p��  �+���w�u�m�:J�����ވ�(�Nٵ��ո{�nll�w�  0����XYY��陮S8����~��]''IReY������Ɛ  �f�  �q9����TU��]���,,,���E��]�����w�n<z�(ڶ�:  �9i����r?�]�p5Mw�މ;w�|���<�������{��  ��΀;   c���~GUU��4�t�-��cǎ�ٳ��x�ʲ����������s  �#�(zq�ر8v�XdY�u�����y�F��]�M�t#���=`i   �  ���(�jUU�ض�k�hy�X�;w���ߩm�X]}w�ލ��ͮs  �#fjj*�[����H�͌�`0��7o����lo�<�᪪~GD��8   ���   {�(�Ϯ��G��9�u�[\\��^{��g�΃dK���?�{���ʥ2k��h�n���R7��m ðY6��!��YְF�(@b�� !6lll� ;�!�q�H�8 �5���=��<�]揪[��H}o��<�|?Y�����H�t�9O���K3�������T7�   �c���ڵ��l6���K,�7nhgg[1�;~����$I�NQ��x     <w    �ҥi�����1�}��\���^����UGY�<�kwwW{{���W   �%�����7t��]ʲ��8��Á>���(�;~�1�%I�f�ܷ-      w    @U�J����s�Xu<�,���>�4�ڟC��kO��;���U�   pA��4u��]Z[[�1ܦ�bN�裏j2���i��'��ߑ�Wn2     �WN     ����//��BkUg�=���j�;U�8WF��vvv4��   �0ƨ�[���Z�v�qpx�t��u���*�xǯ���gY���|�o    ��B�    p�,����1Ƥ�0���n=��ϩ:ƹ��vww���'�\�q    �3�ZM���ؼ�ߊ��1jooO7n<~���Ƙ`��'��o�t��x     JD�    pn���<�(��t�}|�Y��Z����Yk��r��5������dRu    �t:���T�ۓ1܊�rL�S=��4���}i���s�}����M    ��pU    p��j��w��|�[u�����_�n�����d2������S}<   ��)Mӓm�Z��8�B�����i�T��֎�4��<���h     �	w    �ye�$�����Y%�$�VK>�ªc\h������ޮ�<�:   �i���ܼ�^�m�X��vv���uC��;~�1&�i���(^-��     �`\i    �k�z���(�u�EUg�
x�!���c\
1F�FC���j8T   @	�M������M5+U��4��c�j6����i��/˲�}xx��%G    �4�    B�V�R��?!t��rY��}q������vvvTlu   .�F����mll*I����
*�Bׯ?����S��Z;J��k�<����    P:
�    ���fY�f��7�m�a.���_kkkUǸ�b������x<�:   ���^oM���j���+T#����-moo)�pǯ7Ƅ4M�Qū%��    P>
�    �gee�9EQ��s���rY�i���ȗ�.,�|>������彫:   �c�ZM��״���4M���+���@ׯ?�<?�7��i�n���Iz��d     ,w�    V�^��EQ�\a��,���5=���T�J
!���kooW�ɸ�8   ��d���jW�Z]]�:���t��{T���T����eY������J�    �RPp    \t&M����[�1�:�E�����jW�ʛ�g��������+��   \z�FC�Z[[g[;*W��q�����eُ�y�I��t     ,w    �e�K��ιϮ:�E�$�^�⏒1\&8/b�������`�W��   ��$I�n����u:��� 
!hwwG7n\W�T3�4}�s��$핛    ����5    �RI��SC�BxV�Y.�n����~�1�!E���}���*��U�   .�f�y���Z[u@������S��z����K������K�    @e(�    .�,˾�{�#!�f�Yλ�<繺v�c�6�FC����   �MY�i}}C�����U�N��c=�أ:<�������$I��(�+9     ���    ��jI��L��b����x�!���c�8�tp����=V   8W�1Z]�jccC�Ϊ��(Ώ�|��L�A�T�7Ƅ4M�Q�k$�    �|�j    ��[YYyNQ���䪳�G/y��P�$U��)N������}9窎   T��hhccSkk�JӴ�8�8紵u]�����F�4M���<I���    ��;    ��H��o�~9�𜪳�i���/~I�1P��F�����5�O]�    .�$I��v����N�Su�)b����э��?�k�V�e����_r<     �%
�    �+'M�o����Qu��5�M=�Ћ����E�~�@��{:<<�:   P�f�y���Z[u�i��z���+q    IDATǔ���^o��%I�]ι-9     �w    �UU˲��s��1^��ǫ�]=��/�:h:�h_��U   8�F��^oM�����U�>��h��L���S���4�EQ|��y��     8���|     $�^�?���ι��:K���u�}ϫ:� ƨ�h�~�@�~_!��#   �(MSu�=�����jW��f��nܸ�~���3�4��,˾������    p�Pp    @R���c�9���βL���������%�ޫ�?����&�q�q   �'H�D�nOkkkj�;2�[�8ߊ�Ѝ׵����fXk�[k_����    ���j     �Ȳ쫽�?B��766u�=�V�����up����o�  @5�1�tV�����ծ��UG��sN��[���9��dYk�I�|sQ?Wr<     .,
�     <�M����o�1fU�Y���u�w�󪎁sb2���`_����sU�  ��j�����^oMi�V�-!mooigg[��S�0��ڷz�A����     \R�    ��V�4�y����/�{�n����~�1p��5upp��`�NW�    �N����ں���U�ժ�ܶ�vww��u��
6�Dk��x�XҸ܄     \���<     e���z���{i�Y��j����U�XA��H������B`�    �\�e�������j���ܱ~�@ׯ?��|~�i��7I�/���Ub4     .
�     ܦz���EQ�|�#��R�Z��Gyq�1pAx�5��h4*�Xu$   �cI�����[S��*c�5��g4�������gXk��Z�*��;K�    ���U$     �P�$_c��B��,ge��G}�GS4�+��x���&�I�q   pNX{���S��*kmՑ�S�F�~�qM���c�c^�{��     ���{    ��4M��{��c��0g��>�����c������>�N��  �%K�D��77�w(��B�N��~�1�F�S�0�̒$y�s�{$��W     �!
�     �M-I��
!|E�1�:�i�{�}Z_ߨ:.�<�5����5����  �I��������P��f��nܸ�~���3�1�Z�k����4//     WW�     (�Z��?����z�����{����|�~��fw  �K"I�[J�J��<׍�up��O�l��$y�s�%픛    ����N     ��^�?��g���U��v�j5=�ȋ���K���   �Q�}�M�t�s������B�����{�$���|��%�    �J�
     �����{�Yn�����z�1pE��s}}M&���   �I�4U��S���v�M����^;;����V��s���־�9�G%�     ��    �B�j�W8�~2�pW�Y>�g=�ٺ�:���(N����X1ƪ#  \Ii������բԎ�'����moo�9w�9�ڭ4M�6��Yb<     p�L    �I����BkUgy:�FC/z�#U����p8P���x<R��H   �Z����v�뭩�jQjǥB��ޮ���Tũ�XkƘ7x��Zb<     �4�J    ��4M�5���ZU�y��z���sWT^��P�~_�ဲ;  @I�ͦVW��v�ZYiVX����v��u������Mι��WN    ��    X>�����o�1֫s��ښ����c OB�d29��~p�r
  �Uc�U����jW�^OYV�:�P1F�ƍ������crk�ۼ��(ɗ�     <
�     T��$�O�^cL�c����j5
/8ߦө����f�ê�   �;i��li�tVe��:�p1F���ik��<?�c�������k$��K     nw     ��Ͳ�ι/�1V�<Y_�н��We���y��h��`��h�cՑ   *Q����v���U�ݖ1���psc���u��g���$�-�ܫ%��K     �W�     8?����/y���c%�ٍ1z�V�Ѩ�x�L��'ew�}Ց   ��V�u����z�^u$`������q�������qνF�^y	    �iQp    ��YYYynQo��VE�v��xp����1���P��@��@���H   gf�U��Q��U��U�fUG��č�1I�w:�X���    ����    �9�h4�s���s�S�������<���/�H`��<?)���c���  p[j��VWW��v�nwd��p5�������-E~�9��������f����     ��+`     �s�F�~���/�螦�^��el���B�x<�`0�p8<S9  �l7�������YU�^�:P����v�����(�4+M�w'I���|�%�     @�    ��V��$��6���/�v����A6D��;<<�h4�p8�d2V���H  ��YYYQ�����U�Zm~tTl��������;s�����W�y��%�     ��1     .�,�>:���ι�.����[�~�s}pn���>55�ϫ�  .�4M��?:|sp��vvv���-�ܙf�i�gƘWE�%�     K@�    �*M�O��6��#�<�{�����"� έ�|~��}<)�Pu$  pc�j�NJ��f��H������vvv��������ڢ(�SR<     �D�    ��,���������=�~u��E�.��&���v���UG  �X�VS�����U��%IRu$�\��\;;[���;�J�7���(�w�     T��;     ��q����s_�lJ��S9�4�4�4��yՑ  @���'[���[ځg0�j{{K�1�i�v     .
�     \2Y�}t���rνL%��7��{����FY#�Ke>�އ��r�U	  ,�1F�fS�vG�NG�V[�p�x&��X[[[g����{��_�����     �\e    ����j�����$�x��?B�zֳ�\Z�����>�d2Q��H  ��VV��t:j��j�;��V	�0�Á���4���:*�i�k��<��2�    ��;     �\�V{q�g�����tt��S�ee�.��O6�Sx �b����t:ǥ���4�:p��ݸq]�����b�$������_��     �O�    �"���s��{�Y1�3_ȲL��s�VW�e�����Ӊ��F���Ӊb�U� ��k4j��j�����N�tB��������<?�,cLL�䏓$�2��     \�    �z��$�τ>7�h�:��[�s��\�?��4�L4�4�)� �$�Ɗ:�������^��;��ٖs�L��1!I��{����$     w     ���,�~�9��㙚<�Zmn^��w��$)+pe�tx8=.��5��彯:  ^��P��V��Q�ݡ��ĹB������>���o��]���K�+%      �P(�    ��$I~$���c���J�D��״�y���@�b��N��L�ǅ���?�FL  .;k�ZM�Zm5�-�Z->�	�l>�ikkK�g�"cL���?/��%��I     ."
�     �z�e?���c�,��1Z[[�]wݥFc��| n1��lw��*���H  T�V���j��j��j��h�n��0�N��uC�A�̳�13k�۽�����=     �踪     �,��j����B��VWWu����t:ed�!�y��d��t��d����3o� �2ƨ�lof?*��B���mook<�y��vd��Q���K
gO     .
�     �Cʲ�5���!<���VVV��yMkk�֖��B���T��T��D��Hι�c p*I���l�ُ
��N	,G�Q�޾��lv�y��}k�:��"�Od    ����     �Q�V���;�^t�YY��ڵ�����$Iʈ�6��3M&��M�ٌ-� �s��h��[����zՑ�+�(
���hoo��JZkM��[�<���    �K��;     �mY�}B��ǝs/��+X�hccC׮ݥZ�VRB w�������t�<ϫ� �b�,��JS�fS�fK�V�B���������R>�����:��;Ϟ     \�    ����x��{��1F{�Y�u�=]�v�Z�VY�RQ�N�ǅ��һ���X �K"MS5�-5�͓R{�eU� i4j{{[���̳�11I�?�־&��?/!     �B(�    ���̲�ǝs��1�g�l6u��]���d�-��b6�i:���pz�B�: ��K�����7��|sp��tp����m�f�3�3��$I~�9�咶�<     \I�)     eh%I�c!�W�g���677��yMiz��<�(���>�N5�L佫: �"I���Xy�f�F�̿X��(������9w��ᬵk�۝so�4?{B     p�Qp     e�Y�}�����u�a�jmmM׮ݥFc��| h6�ݲ��P��Sy龜 (Y�$O�̾��T�^�:��0�L���������Yk���?�{���     w     � �z����qν��y�NG׮ݥ��n� ,I��:<�Yx?*��y^u, �m��jj4V��r�A��hb��������tZ�Lk�_fY�����ߔ2     ��    �B�j��~�{��1F{�y�z]��״���$Iʈ`ɼ�O)��f�R�� N�Z�F��2;�o�s�vww�����(�<��$�ck�W�y�_K�     �(�    �e�Ȳ�'�s_c��:�Z���mn^S��(#�
�5��5���g�C�f3�����S�յ�rTf�Yh���2��F�e0�N�������R>@h���4���(�^���     |x\�     �V��j?��{]�S��f���ͻ���F1�dnߧ��I�}6�)�)��3I����P��P����JS֞�Ku �3!���lk2��2�Z۷���s�{%�R�     ���    ���j��!��s�Ee�˲L��״���4M�	��r�ox����g���"�: ,]�VS�~Tb�����P���p��f3���jO��RfZk�������2     �Qp     ���jBx����c�g^)j�Q����Ʀ:�R��� nn|�u��lv��|�c�� �Ԓ$Q�^W�VW�V{�fv6�WK�Q��P;;��F��4Ƅ$I��Z�Uy�����      �D�     �'�I��`���C�26�Mmn^S��F���n������lv�윫: H:������O~��i E���]���(�Rfc�i����(�NҠ��      gD�     �G6˲�y�#���2&I���umn^S�^/c$�K�{����<��{_u< �P�������͟k������'������p8(�i��[��uνY_s     ���    �s-M�O����KUҵ�v����Mu�=Jd >,��|��<?~��<��9��c�Q�e�׏J�G[ُ~���J��� �9���������|^�LcLL��=�^�{g)C     �;�     ࢸ+I�7��8�X�
�,˴�����M�j�2F�BB��[��G?=�l.�4MU�Վ7�뵓B;�p��D�����B(e�1f�$��8�����K
     �@\]     �Ͳ�u��o!�[��N�����(OA�O����(
E�</g+��H��d�z�eʲ���v e
!h8hgg[�ɤ����-k�?v���$>y     .��    �+˲O�1����Sb�����ZM�Z_�P�ee���us�Q�=?.�?��ι�c����z��T�=����";x�h��L{{����+�_�1!I�?��ιw�2     `ɸ:     .��$I~0���B����u�]��ojuu��� p�B��ߏ��ι�-��=���
�I�(�2�ivK�={B�=�2�� *B�`���ޞ��Qis���Ƙ_����Ai�     *�\     p��j�W:��Bx�ęZ_�����j�ZYc�4��'�?X�w��体sN1ƪ�w�Z�4M���4}R������/t��M�S�����࠴m�d��kc��y��.���    �K��;     ��j��#!�7{�?#Ƙ�5wuuU���v�lp!���I��֟���^���l�G�$Q�$J�TI��R^�`���#�(����s:8���ޞf����c�$I~/I�o���Q�`     �s���     ಳY��.�����54MS��ohccC�z��� p������-�Gx����'>�yYkO��7��Z\����<����b��F����`0(�����-k�[�s�+ɕ6     ���*2     �2�,����>#Ƙ�5��jkccS�^�-� p��r�K�!����7����O�����1�{_����Z+c��$9y�6������t�G��)evJ� �D��\��{���SQ��5��$I�����(�S�`     �s�+�     �*��i��!��
!�]��$I��i}}C�V��� �c1Ɠ�{�7K��/y����ߏ6��,��Z��9�x��O9��Ov;E��e�'I=��1��R�H�&'�n�����f��;�$�`�]�`��_�b���������xT�lk큵�mι�:     ����     ��4M?Y�x�?%�XZ�^ohm��^���   �b��T�:8ؗs���Ƙ�$��$}�s�?�6     ����     p����w�^B�(sp����چz�[t  ��{�~�@��;:<<,u��v/I�_-���%MJ     pQp     x�[����1Ƥ��I���[����Z�vYc   ,�h4��ޮ��b���5��$I����pν���      � w     �����7��6�po���mllhmm]i��9   ��f3�kOEQ�:�Z�e�}�s��%�     �$(�     ܆Z��H����/�1�ʚk�Q����چz����e�   p���P��~���d\�lc�K��]Ƙ�E�R�     \B�     �L����C_B����I�����[S��*c�t   ,��^��@���F��b���O��Xk�(�,)�:     ��.)     ��ݟ$�w�� ��.sp�e��ִ������2G   WV�Q��X{���
��޹���Z��i����l���:     ����     P�z����������-sv��������֕eY��  �+a:���`_�rΕ:��$y�����<��R�     \A�     ��L���B�	!<����u:�Z[[W�ە����  �Ke6�����</}��v+I�wE�ݒF�      pEQp     X�Z��p�����cl�9�Z�v����uu�=�e   �(
������Lƥ�7�̒$��Ƙo/�⽥       
�      K`�$y�1�����c��^�I�D�nW�ޚ:�U��   �R����4c,u�1&$I��Xk$��_)u8      ����      ��J���!�&��ܲ�gY�^oM�^O�V���   ��c�h4<��B(�k�V�$�(�⍒�      ��E�     �:�O��b��B�=�^�kmm]�ޚ�F��  ���`�����/�}�gXk����K�������~       �w     �s M�O�����O�1fe�_YY9�쾦z�^�x   `!�Qj7Ƹ$Iޝ$������)�       �
�      �M��Ƙo��?c,��M��P�����5��lv  ����R����BJ�b�$���V�ܛ%�E     �;G�     ���Ȳ�;��_Bx�"��  �� ���x��R���H��W�<�!IÅ     �3��     p1<+˲7���^�,���^�/�   ��K��I��n�$�h6��!�      �4�     .�Z���1�o�޿<��]��fS�ޚ��ew   �&���p�~���p��Bα�N���4����(޽G�C    IDAT�C      ��     .�4M?]���3��X��Z]�nW�^O�V{G   ��uS{��_X��S$I�ǒ����9      G�     �r0�Z����{�11�t��j5u�=��   ���\j�k��y��r      ���;     ��c�,����y�_���{�e�v{�v{j��2�KM   WYQ���1.�c�O���B?B�I~!     ��u     �ܒ,�^y\v��c��C�4��jW�^O�vG��E  �s�����>�Nv�1&$I��~�9�fIna�     �R�     ����ݭ�j�Zǅ�5eY��c   P���Ӊ���������zR��-���     �s��;     ��TO���$}���E1ƅ�\o6�Z]�ju��f���c   � �{�FÓM�����e��I���1�g��x���     p�Pp     ����_cLuP�VW�{Tvo��2��S   �Q�������1.��R�_�hS��I�v      �=�      �V6˲/�1��{�q1�ڢJ�T��]u�]u:Y�,�(   <���Ӊ���Áf��B�3�I��'��6��/�M�      8F�      R�^�L��7{�?-Ƹ��s�1j6['���Ƣ�  ������I��(���w��n���<�M����     �¢�     ��R��_����'�Vv?>K��Ge�v�-c��  P�<�55�5�BX�y�ډ��������=      �w     pǲ,��$��{�Y!��E�e�U��9��e�"�  �TB�L&���G�N�?�Z;0���1�Mι?\��      �T(�     ଞ�eٷx����=Z�5�f���ծ:������  �d6�i4j8j2Y��vI�Z{��o�4���|�W�>      �w�      P�N��_+�U���c�v��Yk�j����U��S�V[�q   �RA��H��@��Py�/�LcL0��wk�rνI���     ��@�      ��Yk��Z�Z��߈1.�}^����t��t���*k�E	  �t1Fj<i4j<+Ƹ�s�1�$I�c|���$��
     �+��;      �"˲������!ܽ��nnw�tV�nw�l6}$  ��8Wh<k8h0�{��s��c�H�����]ʡ      ��(�     �
�N���%}�����]�i���now�*˲E	  pj!M&���#M�ӥ�k�	���K�]���$}`)      �(�     �jI�V��!��
!|B���C�u:u:��Y���=  ��5�j4���
!,�\c�<I��c~�(���T,�`      �iPp     �����'c��{��!���q�1F+++j�;�tV�n�e��  �b��\��D��X��@E��^y���H���%�dQ�^��      �3�.      γN�e_c|E�e!��e�$����qὣFc)� �K�(
�F#��G�<ϗv���?���ι�t���     �;@�      F�e/!|U��C�hI׷�4=)���5�e  .8��q�}��h��|��㣵v�Z�.I?�{�2      N��;      .�V�e_v���cC�e������I��l.�h  p�9�4�N4�5�4�N�z�-[���s�'$�       (w      \
Y�}\�u�>#�pO��.��[6��U��� ���(��2�d2�l���2�k��%��$I~:���-5       � �     p%�z�oy�_B�����<���VK�fK�p) ���(
M&cM&M&�oh�$k��Z��1���%I��C       �]5      \�Y�}I��!��	!�.�pk�Z��Z���%k��`  �B�Q�����~Tf_��vI2�̓$�sI���II�K      ,w      \9�Z��������!����e�o�U��T��>��nm��  �I���lg�h:�(����g��+k��%I�����/�      �w      \yY��,���>�����������{��V��Xf  ��<�k<���pz���
Ƙ`�ٲ��Q��g���')V      8(�      O��i���_!�S�(�KR�fj6����[�v�1  �b�:<<<��>�䜫$�1&c����J������HZ��x      ����      |x�,�^c�{!���6T�u5c�q�uRxϲl�1  ���8)�O&G[�c�l)z���Xk����W�<�MIմ�     ���;      pg�z��9��W�^c|v�%)�25���-�G��&UD �2G�٧�L��N�J�y�W�Z�g��/Ƙ�,��$V      �H(�      g�����!|Q�Cϫ��.I�Z]�vK++͓���p p9�5��5�Nux8=y!T���1�Ƙ?������,iVY       ����      P��V��<�������Uޭ�ZY���������zUq  �m1F�f������P1�Jsc�1�F�$h���<������P      �%B�      X�$M�O�1~Q��Sb�/�1V�0O�D���I��l��hT	 pŝ���7c�$I�o�yW�$�:�����j[�      �%F�      X�z����H���KB�Ug�� X��(4��5�L�U�]���k�3���1��y��ת3      W	w      �z�Y�����c���G�mա�$9)���WT�7d� �'ƨ<?��~�q���Ƙh��5��i��C�*����K���Y����֡�Ǉ؎cl�r�#���� � ��5��E��$� �	�(;B6 $�G&�$���N�â�zz�3��=��{溤R�of������w�=    <�|    �L���7z��Z{u�_��ʡ�J��Z���v�Or||�+W�t:=�h �f��b����YNO���I2û�0�gkퟆa���b�I6��    �F�    �����[��?���gz�C�7��srr%'''�����c�1Y,9==���iNOOsz�n���Ǻ�n;�φa��$�]���I�ơ�    ޟ�    .�a:�����I~{����Cu�09>>����n��INN�3��= wh�^���ggg���,�Xo��0o�����'���j��$��s    ��    ���t����?i��:���8^9�P7�L&���8��ǹre��}�,�x�l6�,�����,���f�Zz��j��Zk?�L&����W���&y��s    ��    �oO�f�o%����W�q|�b��$��<GG������q���3�N=�}c�Ze�8;�������e�Zz�[j��[k?��ߒ|o�^'���    �x�   ����t:�v�������ӽ�١����d����]�~m��|~t�� J�g�Z�]��}��z���Z[�c���wW���$���    ��;    �$���f�K��}o�_w}||�a�z<���r��b��bq-d_,β\���~�M6��E��=    pXw    �V��翷�l��Z��q_���\��o��>��3�oχa8�x w�����~��r�����6�EƱ�6���axw����u��|ǿN���    �)�A    P��d2y����$����R�������#���f�e>?��z����w��[��Y.�Y.Y,�mf_�V�����'Z�/����8�L��\.�.�١g    .�;    �Q�������v��{�q<�T�t:}O��?��f���z���>^�����6�˳�����!϶���|��|��|��<=Ғw8    pIM=     p轿'��ﭵ���/U�����\�z�=�m���3��2�ͮ�ߏ����i�Nx�޳Z-�Z��Z����V����n縵�Rk�lky%�7�1��{���    ���    ���V[�[k���'���`�f��6|�^��c��l��|���[�p�V��׫,���V��6����j�:�wŬ�<�Z^l-��{~+��c>�{R�{4    p��i
    p��*h�l�/�����V�a8�?��v��ǳL�޶�{����z��r�د�¾��~Y�ݩ�]��+�勽�$��<&d    
�I	    PƝl|O�Q�[�8�Y,βX���1��L��]�>�t:�t:����V���p�}���l΃��zu~|��������0����\�/'�z�ym�    (L�    �w�M�7�/����齟Ƿ�g����}��m�_;�sٍ���.��W�k�=(�Z�����r�����z��zO��?     p    .����/�ﭵ�"~��bzz��O&�i��I&������i&�kǢx>.�8�oX�^�or�9��7�����w�t���|&�˽�+I�1�y�6v    �>#p    �Kw��O��og��d��d�����d��Z�~��0\;���{�f��8n�^oΏ����^ֻ�mC����ڇђ��"�gZ�g�|����{~����   ���    x��.f�!I� �f�q��r��r���-zv���z{>�p�p~������[�a=������l�{�8n2�=�8��qw��8���<F�x�?���o烙��GZ˧Z�sI^�=_J�����3�    $�    ���Ż7���Σ�1���}0}�m#�v���o#��c���ǹ.��G��*��[��Ǳ���_[�o��F�(}�}l?m�#���oC���5y��$���hky��|:ɋ��I^�=_�=�v    �;"p    � n���}�Ν<�;���?�xnf�ZNZ�I�i-�'y)�˽�q̋��     w��    �.�ӈ���}���iky��<�����\�y>��I>�۾�	�:    �=#p    8����s�>�����8�C����d�������?����1�%i�u    �R�     E�I�l�����1��Z�eղݴ~�ZJ���x�'�<�{^L�b��{�gzϕ�k�k    ���    \r4^�E�fk��q|$�CI�{����4۾��Z[�֖IN�\���$?�b������_N�B�������Ǔm�.X    ��	�    0���!ɟ��)'I��N�/���8�϶֞N�T���$�&y���p��J��$���,ɤ�>|L_
�Z�lZk�$�$������;I�N���[I�����a�k�����������������0��$~��$     
�    p;�I^_�ׯ�?���|��8����d����8����'�a���eȟ��y���aw�l��n����E�=�:ۍ����Y�A�r���n�yk��8���~��jk��V��N&�7�śI�ڇ��     ���    p/��\.�J��7�s��|�?��$�$��f�O�ޏ'�ɧ�d�^?1���q����I&��z�a����I����6��=Ī��i��&o���������i���������6�u���xu:������$��j��$�$Y&���7>��1�z��H�    �;%p    �~������j����(�N����.Ì     �a�խ           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %���b�  PIDAT          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;           %�          (A�          @	w           J�          P��          ��           � p          ��;  ��ν�6A\A��������sU�w �G        ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�    �r�     �K�x    N=�      pw    ��}{ /�� 3s�     �.�;    p����= f�k{      ��    �)���= Ə     ���'    ��s�k�S�w    ���    p�9�5|l��yn     `��'    ��m{ /q� 3�=     �]w    �����<��2�    ���    ��� p����    ����V�i\�    IEND�B`�PK
     ���Z	�\  \  /   images/ead4476f-8cca-47ed-b51a-2c979a8b5414.png�PNG

   IHDR   d   V   9P3�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��x]U��wޏ&mҼhi�������,
Tp|���Ђ���
tF[�UGy�Q??+ �X��2��(�Rli��>�<�4�&��&�~{�u�'����ܦq����߽9w�}�^���^k�O��8������g�;f*++Mu�s���f���K+����N���	�������͝���S���Y��������}����P����޺�c�j�=��ȑ�MMMM���g�V|�_��={LCC�)((��4��  ��\e��cf���f��W �����w�~ۊ%�\�䬂Srs�2rrrLff�-r�Ɉm*GX�#�800P#�������==�����_�ʗ^ikk}J�aۙg����i�������?�0'�z��_k}d���?d����vtv��y�-\z�%��#� ��k���l�P(d��z�ѣ=vf���>E�0�L�H>���$dL*)�R����;���f��=�_���X'�H]����'�~�
��4�	��	��6m�ijj4�w���Sn\���kKJK��L@�1]]]�����min1����	����m�)*.6�'O6��Yf&L� @���L�z���3o;t����ھ������WT���O�Č) 09''W�m�������/�d��´rB��:�o�>D�H�H	�("����l3[-@0��������2����KS�N������ȳֈdv F�L�~$02cEc�JE�����n��{�`хwUVV�A"���#��k͞�{L���n؃�RPPhjf̐5k�)))���;����ޱ}��n��-���g�U�H�XI˘ �n_���f��w��%�x��o?���:���6�m�V����UE���.�����v�3s�i����0�#ӧW��}j�o�j�HZ�	5�w@XT�5?|�Q?Mg�����L��f�� o��g��ϯ�:'�� ;wl���ܹs͛���v����f۶��
WK�?�U�+ ��v�x���o6���G߹p�����H���M�O|Q>��>�V��2R���1/���uv�s�s?��,�R��62Rr� Q0>����Oo�嬷�u�ھ�u�i�K&4��L�\�ӳ���*�_����a?�fr�5��5e1"�}��{�Pʏ�L0VoP� �#�Xv�r���yV�^��M/����1x�'��~�����a-,:L_ �#�zz���3_%�@����	J������̆��g�D�^x��b�����8;;����� �����"�>EMf��bIY`1�Sp WJ����U�餴B'{D����?���RQSw#0�w����x�6������ttt���u�3?3ө,�e��)�����  P0%�zgg�H�y��y�:s:AI �T��9bBʂ}޹��>�����]TTlU]KKK��"%��2ó#�N2*u��ѳ�vuu[�@mQp����Gh��'e���cOW�%m����bjoo�8��E�Ěʣ��6�I�������P3a$m�31LU�W}�U�� 5HݣG;�b���ĉ���<L�Õ�u�<�p:c_i�A´�����++��-�zg��׷mG�{U��}�9ڄA^G�`\NN���*KUF�vk	L���Q]��Z�T"�x6���#	:M�X+�M�z2j@��Y�L������p���~�G�����b׿�>QZZj�*��@az���JB�0`�:��� �ָYqq��I��� ����g �³x&�:�Ȗ@I�������J5�`44j@�)u�X٢/��[�{���CB=0V���h�� B[[�=��"~�E��"�K�^L��Px.��4��2@���R�4f��.�g�9a�Q�,��,ZD����ʪ�0��T�13��
:F���]��ʎ9���٨��,UY>��iUV(4`��@0���� k��;�d�<bj�z#P_�������h[�0U 0����<��_�^��e0n����0x�Z[10�������	�a �P��1첃N��t����!��X7�$C��0 ��UG_��wZ&��Rw�Jk�4*@�y矿�mЛKJK�`��x3�hG��yXW�p����!�D��u�:�^J��\��=W%s�ȑ� 6�
8 ��0&�0�7�~���E�g

�{��
�L�4i�y�џO�tɻ>#	�ݻ'n}f!���bR,�`�x��b�׏��R�-� ĻW5�]���,�[��@
�i���:��M�����*�m�U}񤱪�3u����Ν;��� j2U�+e@��%֕�*a�a�x6�ӯ]F) ���
ߙ�,�*m�G�>�B��,� �B]�T]�`zGG�� 0!XS�]�� p�>��x�K�t�TTT\%�w11��T(%@c������~���p�8���D�Fj�������Z[0���Et!VR�V�Y0F�a�
~�=�5���a:�P�$�/�]K�x&`�HSW?q/R�L�⏽����r�?^��(%@�ӧW3K�!ұ �o<^����3�3���.��3�n!U0Tmq�.\`t�ݩ���o�p CC,����kH'�������u���n��|� �~�`�M@�~-��c�y�H)%@`3N֐��о�{�� �7����I�aV*���r~I�5eic` �YR���a�k�
m�
��N~CB��M�ę�=V��Ŭh���{���z)߾��3�9��+��o5-��օs����sV��3]U���7�F�[$c� �Fv	�����>�m�6��� �:XpXVD���R�m�		��Zx�}�6���R�F��d)��@�����
t3���$��d@0"j��&�5t��d�`�LW�5�Ѫ� AS�x�ֈh4YO?)H��0�Ve  ��'�t�\zZ
{ӯJy.\6��%�x��I�o� �)��[!��lg�M�h��I���V�
s�����#����mI����y�g;U�fr�V��+}��j^�[�����ʭԇcZL���!-�� �q��n)���6��O�9R{>����E�+.�)1�u�r^�JTaL=�������;�f��\繺F`�2�4�Ť�5��!�n˸����s��OL�Ռɀ c��K�b}���_j%/ �K��I�X�^n����nP���Q��czj���1CFWQa��������PSS�y��6���U�~B%b��'��s�kD��Z��Y@�J�!�`rR�v�؉d�_.�B~��
�Mf`@E�=@G�q�u ���c?CC�0Du���G�h���[k��7���9s�Yv�M��.7�Y�ܼ���!�Ҿ�|�n���J�O��lJ��Ժ�!;� R+��gFH�b�J�@fK�c�- ��%��Ӎ�hX�D�o��QQТkRd�WVU��k�m�WW�.�djؽZ~[���﮼�444���B]#X; �c�R	�65^����x��:1�&S�R~ ˥��~|M�C���H��;/�͂�c��7o���^r�u]��l�믿�̘9+ah�2c�,[w��ع�m�z��w߳bַ�:� щ�:��J!E��?!e��")˹󽾛X�Ii�M�c|�d縇�WW��&��]�j� ��/��9��:I�իWELm%���Qb�g���ct��O*��@�I\ E7���q.�һ�j��F*�z��@������P�~oV�D����=���xcQ%�T@��A�#����Ar��zC�ѽ���ό������cx��s�� �L��	9��������(�'�W !a�+%�J����Z���ƈz�cu@��Cg���.���%�������Ӈ���ᦦ�ߢkI�'8,��}��0�!�Z��Q�C�Z_�� �)7x.�eܚ�q\������XNnN`��;���Vk&�x�o���@co������ݷƜ޸qc��D�^+/�{(/h^1�d�����W����3}u~	 �]e�*�D�{�7�������NO{�H�r]�堵�{�5�^��L�6-��*~���{������;���A�{���{=HrbI�+bbqP���YK��$݌�����/NVP'�	 ߽��Ƅ(a��7޽�{�s淐����͟Yn�|k�������A��d�0�C]?ѦFx�J}�Y>s܎(r" �i�h���C�;�s�oI�����)�B!C�j������0���?���~�'\�5<f"�]g_~�eq��0�]���Ŧ�����òf�����@0 ڏnx"y�xZnnN�O�3ށ�&�a2f����8M��'�ta���K�mn#�I�B�� :ɧ2^� 	  I�G��Y�Rq`��;�0�W���eu%8,J[.nhP5G8^�k;^�t,A���ٛO�ſlO�E����pa��#82���}1 �X�y�_"�5&�k{7� F`
�8�D�AEG��{v\ׯ趲nH��	�d�@r�%;���.�%��DI��#CL�x>>�+\�*h���2�&���L��	y�ښ�J�����^q$�����m�LH�R�q�w��lJ�ˈH�n+�-bwݿM����i�HqL��DxŸ�{BJvǐ�S���w����F��am�0�ٯ����pC��6AE@@w��DR`P���h$C��;i=�7�t�[' O����v�/����&h�K�q{J���6"JuO�m��3)�OTQw���U������V+{zډ�=o����n��Mw\ !e�W��W�D
$B�\苮1�^� Ж�1~�_ 挔�����c��� ��t%D����v�K<�5)Q���& �8o��YMݵ����[E3�a�X3N4����X�t�G�
�w]c��<���K�I��[J�0{`�<�Ey(zr~��,�0&9� ��+���2?J��Oq�ۅ��4A-�hpp`�\�>oFL��@2�)H
�2T�W�o����Nzuo�~��I���H)%@t�	V/�|-Q}��=j���2� �1�h$�_ToR��R͔��>9{4ka��Fb\*i�4.��j`�4��A��i"MȦ������~ƕ�aRK�J��䏌S[��gv�d=��@pY �#�r�Z-(0��=����I�K�.�Y[�I���\t�֡Ȯ���{5�bMq�#����91��G� ��;H��&�Əm='C)�٨�D'R�l���#]T5D��a~�J������䬱ΰ��a�G��0I3��IZ�&M�,�B4��o���Ê�ԍ�C��s'�?�7o���^{Ռ�F}`'Lߔ�KZ&$����,v���à�o73C�#���|
RB; Oeف�t�����o�J�����ˌ$�)��0���B"G��݃�8�s�>�	s�	����,��.�sRDRԱ�6�b��P��l�Y�E��{>$�%���yT$S�'�g{�����͠��*k2�����~�ܝ�K5�]iT��--��h񇥜:�}.�r�� ��)�w�u�><��hzhJt��K�	�yZ�@ϣ�#�é�g$i@ Qi��޽�Tiԧp�6.��)'s��l7�$��UH��Lti���Ž7b�&�,b�c�!5 �=��u�a���K"ɠ��@��fs��/�r��� �nFK��+%����r�p�1�5$B8��Ӿi�$'�Y��U8��9�钼uo"�.๗�D}HC'����ʆ;��5]����-]z�kW��'iy���#�qΖ2#�{�X2��N� �w��:Rl�a={������ �q��-�@�7m��
��;M25�ʽ�}���>}���qr�Ai}�L�q���'���BϠ %�w�Wa���T�:j��}YH�n2���~	 9I��3�L^�~WJo]]��P#��䭗��:Rai!��)�r��"��P�S��~�z��#�l���k G��}1R�9�No�%�LThM�L2dCC�'����۲�V��I��RJ���|i=d�`�$�����^`V>,��b�۽ޙ�<���5�ܽD$���.OMդ���̈,⍍�����y�ס���(�o���5a
��Ց����"�����ވS肉�m �{�_�'��'�/����\$0�:w�;�}vc$B�n:n/���6)8w�҆ZX�Q�~Bl��7��;�PK��$K<k��iv�����[�8c�]�����ģ�z��]RI�WJ�I�4y��󚹐�N��y��/O���8~7TWW�{��W0�1$���Q��8�IG�nAO�{�Y��M��������uu���<�-[^��4O������s���[j���f�_�KҐBYk�������r�6k�|cL^�>&����
�<nܺ2�����Ps�X�{&�zݔ�UD���6�:v>�t�^�~Æ'齹瞻�nMţ1��A�08���i�$B�\��R�0��m����{�Uzf&*�H1(޹Z_�7�imm]��ԸZ��������u���}4cH~KGJ��+R�koo�IT�52[�8��ɩY(�>+}� %sA=u�2�W|b��[`"������N�} ��M+&��� :!�a'�Ɓ���/���XUVVvEQ�ĥ�;�����E��w,�67�ąPb�p5d��z[����ċ��S_?{��#���iv�ޕ0�{���*�pq��Y�p�y�G���oϞ�� �j�\f��=��)w/��Ix�h�ß��]�5��__�H�fb�0�I��-��:��6g���v�4���TOAt��K�Z.?��O�Đ0�gqq���-K�^{�ʕ+*�[����YY��#��_�E��Ͱ���J_a(�9����T�N5�h
����Yi:;jW�������x���?�}8�`@'/�=��^�j�o���i����}�[�Q�#R��wn5�2An��\צ�yy�_&��9�t��X#��q���N�'��~�0�KԎM1|B����������á?��/��$I���᷺d��`�K���d��I@��d��I@��d��I@��d��I@��d��I@���stD�Lr�    IEND�B`�PK 
     ���Zf��g  �g                   cirkitFile.jsonPK 
     ���Z                        �g  jsons/PK 
     ���Z^8�H  H               h  jsons/user_defined.jsonPK 
     ���Z                        ~{  images/PK 
     ���ZP��/ǽ  ǽ  /             �{  images/0b351edc-7875-4477-b820-546ce15be531.pngPK 
     ���Z$7h�!  �!  /             �9 images/e0155ecf-753f-4e63-a512-9d8bb2c3e0aa.pngPK 
     ���Z�j�7q 7q /             �[ images/b909fea3-6005-4c04-81af-b407c7630414.pngPK 
     ���Z	�\  \  /             y� images/ead4476f-8cca-47ed-b51a-2c979a8b5414.pngPK      _  "�   